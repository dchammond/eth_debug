`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
L7mrIa9gV/8yw38IOlt2y7xFlP71OWjo8fN/HsvvfP2uXQqADJ1GDR6P6KJdyoyi9pw7QREy+/bb
ykHHlqlVOg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
txNNcsstWATxcfBvD6w/d/CBhO5fZjcRz/FaqVIPXI4mHIprXtlq7mVp1J/E109Rnayr7yVNWF7+
ovPpXJsXNVhefw+5DiN2s+0nwS6xSE45Ag6EjmROy1BmSx0nLGSNAYFmNxdMUxU4nJKCNdkpqP2/
aATfZh4/1/ULWEK7/JI=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NJe0hXHep5jeuBn7cRVT+YGR8eUF1xQ0orT38woIC1xz0Y0lgowxb0lNuAdNTvQAntxu3uWXRUo6
1UeuuzrWaaJYwHk0iP2XRBJdtm20A038cEZQJMEkAGZJFu8x3xTtV/kXgd2rVjKyWxt9jjiY3yrt
BVWUdwhCCMRHQkyAO6WPYA0NNcm6cH1eztOWhg8Qzwk/WOrBHQbL99RRhAdkfTDOG1ZtxtrWoWGQ
UbnAV1I9qc/QE0AExKGOFDj4qlcv6aoE8jBsgfu6DXXXGO0FFAFgy4vHBzg7x3YAu1cIwMcNDCrA
cB5dATMd++vcmJrsIsTKDGq3429+ZVhDJuE5gQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fH0EPjz2TYOzRKzbqVvOK8tpxEbZvVhUQf5CDZAfQEcZy7U2klW8EzJzs8E04vEa5JNwLCByhcCH
WR5dbm7D6EBjFNcp0iKrCwDVQ9UmpbECY0n8OyZ1GaxIEIxBmHTiYXT6cv6q9LCfymLoa2t4KIUP
53Io+5as1cH01bnS0a/c3xLrbEK4SaL3kIVQWOP9dsfF6S5uHzonbNt1tZq0TBogn7yfO0DcJiqY
Vh5ZwyJLD6OgKcgt6YyEc9CPEo2Cictg7PzZyeA3knJhGZzVObXe8tKAjJqoM5ef+q4ZH1f26z9q
7iHSmXYhYliLm3D2/pDu+gSENefhG9lmF6j4TA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
oKosXxtRcrsJw4OmFZtAFBEiJNxeuxyG3ZsGYXF5P41XVqq0IHrv+VhGM/QALKzaS1dhEa8vUfb/
GUYGS72iH5U9M8OJv9BH7p0R5kZD/ZVD/OJtVqnYYmQNajLr4P3PsdoNfYfgBkqfA47gfpapIXiM
sTZVKfh817zbsOdsLBw=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
O/DSm2QgSi+o8guVg/zvFTMk7+x+wYMydsyZmhosYYrfaE4YDrlMnpcNPCFNgB3xI9WQlGdy5ZcU
fyzIPCgMiNfEW+skbXWXdOPQVUpayFwEbYcrFylRjBtDllOkTO0rjU0wll7RmdQXLQUzT+fYwkka
zN6jD5ApRxkk42jmRTWsY4An51Tetw35MbULnzNhq8bw9yMXzWe9KLIy2VDC1hqSj6V1aDMQjuPu
BV0HVYNHosBJWNg+tyFYW0bC9b1+X2FefvVNHGTFaRBGIdJ3SW1LOgWyCtR8uD/SWEKk1p4Oa++0
Vm0xzQHxa/aNBa6tWrTOY8gIkqOSkVLasM2vmg==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QqXZjpXIW6Gl51ZwyEfg2tycetjqR8sjVKEOc9Ie0VBR0pC1t/Yt+IXrkkCJ1qs945fqBsTnRX+3
n1xf7GqUGzuDCeB5tCUjrJuswY0bBDGkklt8oRyvyvqYu2/P42wbhs5NCkUhFe2qjMS+hCqxa0Rs
RpfbmLIVcBkrbn9AKX6G6ayAyhalnq61r0rVx3ttuNtUeE7auSBcmZ9gdUWbqgCjPPDTxXC0oFyZ
OC1MX7DQIJ011ERSJSXJDjUR763YZpPfVe4v86jfejPELIQ/mTVE/qeqyldz/fJyaAgbjwjVo9+C
Eua67xq/4bYRagYL1IkzMna37u9xZTwbs20QiQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_11", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SQTfQj3cbELfHutu0HrpwkMbEvVG1qBxr0ynie4656Ymvhd57Ec/aa9HftrkF/k707zPWnMYYtdP
EkDPJVP0CW5H/v+QOPM7YtEHyVjslb/96ahBvioJ395xBXS2mo0kuxk98xOh6BHRp1rNGx0d5tz1
wXFVqtPvmGXZTdKJgNATqZ7huJpWjU5XbVvkYw2LxNJN47xzUd3rdaLWLPPu8SThDlGKUzioG2Cd
oGQYiDNCFuuNmtuHXXWi3WV2PPYh3oCOyCPNv79gQRkjOxggSz0U9xf/BGZp4GRWQg/AvCLk1oPH
lkt7yxmR6ZJk8t4k7nQFLt1s5Pm2P18xbRNloA==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iIA4CVL/b+CBX40HI+oesJIUPmd0E1IINOh+7nGwlfqK60HzphgoQ/rhA5ybsl9uuU4DF1yUlFgp
qRw3klLWCRF2LNux2TsySGaGpqnaYrVJBH0FSz7329pSDTljFKOAU2jXGnh+15R9zZ/a8Qj1SD17
Bk+aTOax62Jsvf/+OyD5a6ga5tMa7mF1SaR8A//+oqbfJ5iFZKl2aGQnNgXhVbw7ABA3iADvXgop
zbLtP0BZ0EN3jKNXwv1Cw/n3BVhfmUYpQKC6Tb5YW4DO+vVunbQWxZi3kKwFfm/oqKU1Vy98wCJ5
J5i8oNRIzw9Fa+oaHMI0329PpiKuT+LHmyBzjA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 860576)
`protect data_block
Y2/hzls35MdSmztEEX5tiunAw/9xht2i/Zchf2xmso42R1Zp2xM5CE9uXikoFdyVxERvsEPtZTiw
21RdhmA+2/J8p31Vzgrd39MNg6lTr85q4pd6XHXORr796OzFalkkMQte3frr7IHB/ZfZIQ54JhMl
EwnVLyoWCk8pFL8JywlZJRkm/ZTpOtMPxsmE+BZjCGDmIdKTBgSGIZKmFgZaQd8AIHdg8/LjVHcJ
xpoMPdPidrIPIuTx+01l5mJ3A612w2SQoZQ2QwhXk1n4R5zF/uUJ5Pv3Ex/qzio9iLFHlVlCM17x
TgoEM8iyhl5k3Ne9MO3qNQylgBXtSUgR8DCEJ/9U7b3dcy7P0NHKpXS/oLizcv0ytkpuLtuWzeqj
HTHP5gEvvJjkgVTZKsOB4RtMdzMh54l7CXdy6o/QJG161FpKg6vjz2sdz62DCobBvIBLI1gHW821
RPiGw08LcfmP1+r7ko2YbcRYjxBzgMy+KZanRBfqFeXqqE6Y1GQLpIn+oZQgj7L0n2lCV402TVkz
kVyWP1C+Wg/GeWwmb5+yrCQ+BTrtQJpRrxEP8Ls67qQuZWJUz9+FJTcL0ycTSiYd6owL+ItLlT9f
S5/DTwt4fSNh2iClQ1k7l8C0PkMGwbtYApgdyFTqloEsBg9OX9/voeqMfTlRxQ3qW2j8N719Dgto
YohkDSys5xGvFXfW6YUSA6VEqZ80ifQ79/NKgIv7Ja8xZcnODw7w3ynfGoeQoYXJdj/4Dbc8FClJ
3AHu+92s/R1MFSLZFLfnAA9UqzMP3F0zi03bkvF7R6EMN8uoGfLlmEHvQ78Wihvi1XBcttyxW//E
R3e8cpMdw2aU1msxdsPbgJvIBlIDox9aFyZUyM0hb5giFcMTTTRS2ajMQfXUEVjvaPFeHBFvQPJw
Ujq+pHCE0q6oDrgkZjPrmYS+vyCB5XPMx4P71auPItJB8DDA6UTRkey0/ZeavgIZ3PBaMZhvCV/G
LH5sIwgka+r07PeIXvOEruC6WC8bvnLxkW1KvGbgAwFAfHtkGZlncSp5qCf8Pxmxo+ooYsSV0L93
16468Q9tAalDrHBbRUvwjINQK+gPFANZtuEMWzw6aNhjX4VMpKKf0efhaG3VGyO+afDtJUmavtVk
LlkaPWMMtBWSpra0Le5nSxo/+7N6Y/i6UONRC1/lO2fkYUUM+si/KxZigFj2zaBRbGtDD3KB6vJd
Mj/3QwlvvX0aAlLOV/fkahDvNtiQ3MKi+qpIQycd95tEPFhyGN0ouDeI/j73NR2HzIKgSGEcEVF+
mQSGNDnx/tU9+7gEj6v7EKLOGKWUNvDT24C4PjUSwn6Ivvz1pH2NMdsmmXAO8XB4M22v6okibX+n
v3936I0IQOJDKjsQTfHwY9CcNl5ElFqzjvbmJrZcOLV05ls/90i46BRCHQbJgu15xBfWqDxQbvay
VlcZMzFcGSgsy3J5+1J06EeadfGcPPtWczSOEnn1A04uBWeDQ/5Ti7BDWwp/23pbmF1FBGF4C+z0
6K0eASOVSzBWrCiGHF1iAfi6YvTBJK0gFEsXRx04SYl1gMkbKi7Tyzu6yQtYjobwgm4Tik+dZNfE
MNaWrD/iqXhuQFLVDqQGOcVYhdPwljV31qP4wQonryxEdDWOYLxbqtPH5IK7ISO3qpV352DTaaYJ
LnDrNe129Sf5WeMF0eqXGIiqZRdnKwsL3hCUOrBSuUcg75RCY05ZchBYuKL98n1XDcRib/83P11f
44iR6nPdnCwwlJcmhwScz1xS92JGqK4B52KK49InxNX7dZ6iyVmkTJpiPmC0VBz88AZblN9o2bVv
AXmzNiwVkIx65BP2e6dUOZ4IIP2ohe/spoUyalvdULotLbhTgT2vFrtDF4iQM43b/m4ab20dCDyo
j7C2rpesAqzEzCxMvOR3zyerC3a7xsma/Xh5rFyD6XJ5wgrCBNdBLZ0YPMuVdvcLwJCNDieSBLsR
insq6SjhYpzIQKLABX3439CzaxmaCzHUtJYBRLe9OAUNcMxjBfL2hims4zV6RUsCBp0gcXEKzcmg
R6sZrgnb0zQ9vZCUDUPctEdIX6lPMs+QcjOmAzXakduzx+pIFzsnA9+utIilF0phOcdXK1RjPqms
bF0G4FfwrX5S5SXlcwPNx5x3NZu3CYSTCrlVRZdLkYCovwmRNYcP69bk9ny+dXHvRJWNQa5xZlCz
7DVBocpVLaFdm7eNJSS/T3M0C75fT0ysBJr8ohz2rKCzDSl1lrxDX0R10+dHmLMyqkKwSSKr4TqB
BOIQYaXbs2sHKyMCwTzMr83lAZHJa78PMs16tmKL5QSpZc2ehfV+hsi1XvX5f1fc9Int9cLW6mYF
jy+FhBbP5WGC6+xmVjWmJBYW2P1lRjRrSRM2dfYd2DbJZBIRLSGI491oVZ9z67ZFZhdplOKuIzVU
I9SdVltPHAz073ER0+zn2zgghH7RvKPxo90PzH4v+lPmfLM9E94zr2M1E5ooKxk6bdp5/RjI9KRB
RbjmN/NS3B92Mg25XqJ/UO0XYeJg6n7fa6gGFqm1NGLiMig4DNObatXlYpcPNs3yJf+nGE0BrTzV
lZyGAkUsabIVvuXKlHhhp+VpMfHkHdNGAQY+byGz14ABRpdvqSqh79ueN7aStQsYzQK8T0/Bo8I4
YjW0YwS7boUiitBdhnVastlo2E0SN2tRrmy5dLdqq7JJ7anPMDIOxAntbRqW53yvLO1vZrmrGuDc
sPI16g8+bEQDQ4gr9Jt5oj7DkajIFbvEsVkSI0pJNOMowBK0XVKwVIJKhB8dik1oC1k9FpMzWunn
4J7Sy4475vJKz1hOcGsxJ2tso0Lguu/htdpwcfOlgT5AuIssgkTtV63+DRE2TJma2RiSxD9svCea
lhgvIyufvG6aSxcifxFD05biwW7HPh4OyDfN5yaMWImLABsERVhgWNlFa+j5o+De3KwNUgYHGYO0
Y/BEKRitx59UTuWUEC0GvoigdUdjos5e+f+/6ChugK2dga8kDZi0rBLy4smH8sOlsd771VO5d+Uw
0LMPUgDuTuf464PQmzr08nwAVGYDqLAYUoBgJRlmvGKpTV+PxxR4BLakOuZ4gFgZelcwnu3lp2Fu
l6Old7bsx2HNDDpMkAyrofBOfS4Kp9lWDsU+Why5f+F/UI/4wwjubO0Fc8JufRO7oLu71K3d+/xR
q6mCZEwHQu78a6AUzXQ0o2qYeO0xpUNd80LNEAQl/BhH2mt0Nq89RqP42QUCo1yu21qlzJYVjsos
ce+IvWdSPOp+de4XLftMqOv0dPyYNfj85J73Y6ukoUNFPzTBGVuBbFfHpPz0JoZ18mUxt9THoI66
LMAONMHBiXDBZsfqe44xI4LBsVnjLYeRF8iXbQjA1VwAhfVp4e4XO1nTe2wkXtmC55G8uUzVvVPC
5B2LcWe5xUjQtRPnreCUr+pSOfoij7TavWaToDdDgzG9e/zflxlEVXR4ZHM+guFx7mvG8Tb6S6wX
6Nsf3Yuuy93kg7oDn+E7lS2ny+yJqYg13utv1rmYo0ilwEB3/zlpTOBfTWC2C9/HgW/95lLhcIQ1
NBZZSJvYQT85BJ/wAi/4WejZOU2iwabne+fv7b5ChtmJzfMM8O1wY+Afn5SNaT8qOfQg1D10RsYO
iJVlxcGpfh7LJjmekMFgWLqgC/NicDeEt4hfLB3JJvXYIiegEoVZJjQIF3/b5t1/keMVqAsHpxnF
OlxrdNQ118Ltlb1LmwhVzA9YqoSRVK+Jgz1Dp5BKnkQjyct4yMPr+2e1mnpm/Eh2NtlJCfAfMt7R
YCyPNlxxq9eIUouB0WWvgdmVCjReaytH7JlsQu4SkVRrzmDD9Kalq9fCg/IPVUARVlqQgu1frMCD
aQWgh90D54Jnk1efnE2XeHrTUQuRJOBL8lccp8BKAIxEhk+VC59Rw39YhdEjdmuMSDZi/J2MaJ/h
XMDZ92DLx/KGehAebLkCiQIW37n47GA5dzMXCP1ZbJKCmJXuZaPYgtK5CUGnS742TXivL2Es8U2L
pi8Q9ArmFrMkYrPHY6QbSCkKE24e/JUUa6SQcOOfzSs8/fAPH/O9eVXsFQbC/jrATcgdv3z9jUiJ
i1P2DShKnimldNhgk3QgqVD1fSCgH34MWBbdKVit71i7NTr4NzV39dW7ZDQ0Nx3b2EHHM/FLptR8
FuLEuK0hU96XCI8YVu1I92mUwbUEmKGMLseIF7grghf2FdH+VNQjpbQ3n6Md6uVya0dUHpRF55Ct
J4SL3QbrXgKuRjmXeOu2HJtMQbozqDyWlNbiGOyCdriKkRRQVU1yxTJ7FYthU/JeX7s9tybekPij
FgLXSrB+CRwzRrmosOzx42zmk7CRrxw/vDSl5gAgSYYoCDlEbGe/Vom6GvASTvlktPJ7uiqGl4/Q
zQ0I+7isY+Tz85kxdS2YEvHR4ARPETXIXuDdn3qfU9vByLbSyTK9QWCax/9MizxsKVNK6MgP0wMM
FhIZ9SeJLmfziXSb3r5xUGJga/eYWlmY3egGLeuO+HeLU/At1s/6fgiYirGXesAk36faPjcbtK0m
7JG6swlZP4Ib1eX10mEii+lEyNR4peDZ8oiSalZ1TVMkiqqK/qU4wtIneW2cBvA1YpQEO0MBix4u
4i0eC3eDl/i/qehIvy4LLNnRtKLqbFnllHkdekMSe8fFsBVR3fYRikNcBO2Jd4ke0EPeLBsZGgcW
Vg5UZEixWLxT+ms6kv4mVqKbM2evHO2rd3pSXFPN+BWskPYt7m10dUyf5Zayte0Tr0d6piP4FO3E
33WYJf4Vc5ASQzHbuEa/QR2SE8wSbAQ0+hszzpu1cpIJmyUvqdfd5IkiU22xN1NPKNIvw9edjYHj
oZGY895dazQl95f6JBg/7CnseU7C27XjhjPrDUg/Z9RLek7GNOsMq44nquJnFLWOhuba/U5V/pIJ
I4LZpol14HE7gikgbP2A+HhuLYbjYqJ4UknFQuEt/n3/D+uT2tA7BmE3zP+P+iWPgh1gtyPhVhfh
CZuTFdS2pqAH1gJMR1oYhQNnxQVCauZ9GrIncn3/MbbcsM+RVSVuUabKZvEQ9FhhWpE23xiSKfzu
bTi8vFQl4JiJ+btNBpXcO/8Klbsn1N/qIcgankvCkZHs1fhI2tdHJFLgsZi0htmJf+udluBBV96k
ToAeAlQ2TQtdTtpTAihh/0IXCWn3ajzwbdJv5eEq2YlflaVeOq1iKMWwmPiQTnC6NkXab8IQcDmH
6rdaWsZwa9Q9fo60ybLZsZ9big+bwv+u25ElDRDTnQWby9m8u5D9FDJwlaWhZKn69oxIwxPn1Fi/
bTfI2gPpK45clhjXhR/I1uyaBv1APbNN/db9nosaX92AGkKxCzYgiFqGI9FIbtjlwb+v5SzhfQOS
Boqbh3cmYksOKY2DDkohuSiw2BGFaq9oc4QfUqguBc7sIA0a2rXzPTDaezUJ+gJHj1hH5W01GQD3
lolnhhFY1QUJLDxBRIJQMhRnZFdhC9ZzWWpt03Xtu2ZKkqa4YjfvvlTVLed/YSHvEBk3Zt9jRow0
w0V4hj8saSmmdyquKx37PQRt3rJsXTsJC+R1w2FZUVuHC4ZTsikGXdG/WTBPUJDrLVz0FuUnHe1U
NVVu9WO2ZIe4uEJsu4Bph0pY0BNwIWPCVlfGFJVRrNhkHCO1556j6FdaBTIpih3w9Bv/Z392h3qz
bpX+AMK9P6lXbVmRMPnpA9qdINCaphamRw4qR+5RORA2otaX1Aaqsnn/F+ZPk/QUH8o5M3DcR4y8
dmBcb7QKKh4foqFq4EbL/aSFnbXybYE+UP3tD6hPyx+x7qmLR5tzoLIK6sxcYv4nxdmO35CD3eVT
00ZqahM5VmDKIwE7tvUTFMcqbV8KzDKre0ZNuSSF3PiMtHFMFzQQMZkBa9HpuB1+FlMClsKt/2jH
M4scasuYUTTn8IScYZ7ZUlHHKCp2dnh/BwA6QVup5U/aco4R4Y4trw8vRoRcyk1mnIUYgitaoa4C
uBH3xhYf68BCdBAG9ow+0/CLqqoJsKm+BZazGtQD5vWr0rc9z/Ff19URZ4jKPS4iN4dSXnmmsIZU
x46qlPkRx/UuE81wiFrDOuosyRtHAZXaXjSfOIo+bNEE15ZQHhbzCzjAMJNofqGDLmFNBtoR7TcU
h/rldM/Yw60RUvGT4T6YFIbAcwDzrCdTUzMAyJtrD/XJyL9QB8cK9fIkdRWZOqOL7WRnV6SCzVP1
l/bZlTB/NXYpzFPlqwTbJKK0CyTAB8U93BMBoeHodK1ZiO5mtXAGc2xjPQglhK4zjIHCqJtIgSdx
XrQAga23pvJgJUcryaP2KFKtt8xDVoFAUYkNFggchQHpXfDewj9+r81P7P4ASaMoyoVtEq56LREs
r83eESPwOXDgwhvd8HCKE/7TBsjDK5QMDEfa/4zJm7WEwDy/Ku4jx+QFFxWpCM2PcrkGQLSCYuJY
R1WWHHGFPLWUMUYXWfqZkxZPGg/gOYCspdQO2RzsfVVVPCnHqSlHmE4FgLk9Ff7Q0jHvFzAqq6SU
XJj93ffBydBQ/m9MAv9oZA7EBVo+m+Hk3+1vtTCtpr81DLyojAm837Tg6xz1FiAVN3eV7974Nsys
2cSj4TAzwWNILh0HD9ju7uL8KQW2baw3SR2GnnjBkuJZCE3MIOcnqzpm7n7Y4sVVpjccDCQafMpW
UGUEaQU0PvZUZhj3A0upyMXtZ5hdGlHrk4QfK9jcP7U+jnf+FBjKwjvsSILLXGdz0CHcfqOVsdb1
lYZf27gvTaHHUE8QTL3XASmx8LIDv+7TRPQX7HhIr1GOBF3N0lFBVPcNU6xjmzK2Gzlj4jAFCeni
IQNnb5puC6dF8HJ9zXnoeJGuYCJGupkCMA59AzxOCZHXPMdf8mvjjlS5WFxUazQGqZjvZaNhF9Rm
gEk3/Ef/kZiIpTh5pqHXJalNd4cXEyCyk76g03JVKp6vzPsDqseaN3An9+dAIvAaiKkDw9t07nqT
c1VB4CK0uCQjrL3uNbIRuS3ttP6gBfP6AyRHAAECs0g7Sf5PLL1KGIbrwVtp4ioiFnk9uYLeOpR5
75nIUiJmdx2/ib98pGOAnGLdF/KXPmGxYXoCCon7x8VGzPvTEl8J1ulshXrHEqbGO0YI78vQDNXf
TuS/GXMSQsIautv1ZxJXDuXvceJonPNszJHuYB9Asejw5UOOEsEx3YBTdJg85JuuNjIxRYKLNpTT
BuhCuj0wOLOuHgMI7jAoebWpgf3DvYF2FkS7UqSgIr4cY055nmmLzPmJ1zljuPXsIF30PWdjWURo
jH85iigFrEnruK0If0oUywc1KhWXJ1/2u7GLWw+2ZOPjJROf/eKjAm0LARkWrTYYx3c9kcHBopM1
zhdxIgNVivn9z7meKzXNMx2psZf227Vdqzgp2VZ3OQ6TW7RUcUIGFGlpnh3lbM8uEeXn88JYVjiz
RMeDAPGnN84dqaO7w+KOX79hZsQHgyU8lEYd9LOP1V6DW3Zf5WfSxbpBHtQNStsyHE/rNTzLQQBT
5MxQ86ciSjQmA9oLiW7sM/8vBOyiD0Ehq67DVvYUzQI08vUEsEJQ4C2NTz9G5gN2a8ZseuPK8rte
rFfMTTRtKx03JBG9a+npz9+RJgkDXSQrlW9o0hG2qMuNbBG7GAl8ckl/z+fvzPLixDkqDzZpW95i
+ODfZ+76VI8dVS0q4+siM9niYMIHB9jNGyCapgHOxwQuap33c7JiT4K4JtVVqQojL5PUBxsM95fj
RDMTucyYp4nJlTUoLbmHiUB8MnFweYinT0Pa8IFPxTor6Wu2SnadPmCt7E5YahSQp6NgHV1AEQga
S0yRfNBO2+swnfgVIGsOGo7ZN2HRcZkEkjmQb2noCrGHiJ8A9fwCsk7nRrT+vdLH7qXcs4iX4PCJ
0jvfhFHfsv44MYVPqG62LFsplc1mB2AcA4lh/u4z4nX5PZeKvAm4anyPXpnQwiBQuv35SK8O1rii
JgOMMIoRrM/b7LSKpaOoi632yRPf2XU/6FVhlpkdF3in8pninbQnYNceeH6H5+G0cp9jbzvLQSP3
enMAgfyFRW0VRC79mXz4ahqB/GvG/0RSBg3gwhGpwdlJtQWvfGxnE276j/GefMEM3hYSIxf8RudJ
c1iGoRAUUpnUts82KqYKwJLNszmcbLI+5P8wazGV93SDW4mdddmrUwjQ1m0e5ZcvEe9ijZoyJLVy
kRuiq7QHR6bDrO/zIDTPEZrj+6AsDgtdm4jDxoqNnKGbeO8ktIXcfDLhbVG6NCTP5yJVJgOrCoa6
7S4tid5lK5KOlMH5D5psZh9ykE4CwRk9/ZVBDejn1Q4/0b/Fsz2lz+uR6/Rw006vkLtMbowDVp1L
6ElsGuFgYFziTx7ZzBq6uJQUKVqO9U3cUSrtUvI+cbHz6buO9VYJ4L6skwBPaeqNGDqbqX7Fgp5H
u/agCULmMJytlcxAndWz3gfmuaR3i+wazDYroh0ydM4mzTnljA12USfuhxmerkUljPbEmNkaBG+I
euQleek0z4FYdComVKwdijg2NbIhZmwsJk5G6pydvgxgpWenGWSS5GiUJJ7rttEn2k19BcVpdrKe
mjOSAP8BMMvjXuSSyqleAZHNsGuJUi0oVsLeOWGySI4d1H21Fpw04FhAf7mH16GhTcTi2rejgeen
H82CSja8LSQmN5FFLetkslYV03yUzN49ZWL8V2LBJV7pFy1zKWRmwsfJygoWb8OjNR3GZxYit9N3
4BzgchwE4pTnFERjuxKrXy4AhNQa+jdv9vd/xt3GSf8gVjBz0rZD5BZIEXK74uElSETjwlS28dXI
w8+2jr5xwtsvcvHKUZsqBfCM63F8Htl5LCgYntm0isyQn7SLH/V0MUWm3x8A1q8ELmwxes9CsGo0
Dmlx0CIQEIFeP4OUb+p7aMpOj9V6BA9WjKKlgcyB08lceLWCDq1SX0aByKKUX/nj7DEXbVsldUBX
OuCvLOF8LlhYwHxZrb5ql59V3wZ8N+6ihB6aKcdBqobBGxsq5vQlEs5l2X8tlOLUrUwB/mSZNbh3
rjYQLDn0lUINCj7m8VlHQXsmjTX7F0hLfa+EpWrmpmH4IZD6wXQAo9M0SqPmjtpHp+VggyE7OeIV
H3Xwi2J9Bw5PHLy1a0cmJXXga5NhnshzYFmG9zXb329uMgQRNefY9R+fBaaLxg/rBEZUhkUBZkoX
Hcb1dtSq9IuPCuwI46fSyvqtL7GdaAwT/vk5N9JtmbQSUNZkfYVDg/3LZDohZX2aCTWtk6r3VWEK
3IPpuP2VV28VEZoMrPjcwUbUVTwzxXHwC4UWzFVz3WoJI5SMRqxHYy0MpF6wxDfZGNxJLKKy3eoq
3iM3xi8hcuuWiNhHa3JM95gDMPdg/Bu5t+zmpusqS3U7UUWpee6r1vkJDjd/f0mypofRyCSWTqS9
3NCg0LxX9mEflqqFQpDTreTfiT269xwQfJhSFweMxZadvaMNpyFRqTINjaysC+AYAEJvbeKP7qCR
iC6O1JNRzHz1PntpRsYhfHvw/ptRFnqFeVc7GuMcF6MWn05WRHO0zKIurgHKedNavkRbWxx2yj4K
QW3C9VaBMqG1H8EOGriE6sFN+AfnqwpFFWPFDm17AyITSx0EpneQIxfLbmhv+/l+bvxDXqLG2QxL
ZghLWEKFMN2m68mMeuSvv7naIDfYvNpqpVZ2c/2H5IV/RrXr4QGwMDk9OpQuejMlfhTAXgN5UeTM
DLRHySybqyZMIm6esQvzzB4UMeioddHaL7xb5PRf0oDSFYHoRKeNebajRmQPHc5YF7Cing84iQaI
FFy5wfUQMEliII/DMQmIvoeFktHqXvN1eVaWuJbS2zDt/ivpRpMN2uzOmL82NxUy4cPnukhG89+9
Fr6ee8YjT1KEFLx+Rdi5cALPf276fujjDWYaNiRNSqti/S2gTIKv3XyU30sUsOD1cnydcIe4X5Pj
NKEzdCuPZ3PwMqe2drHBpKrQyRbAN5RI9aw9/Li6F4vFrC8FcCPuiyrrxkDz5CFQAl0rV6Z5alp+
X5+vsW3Sy0p4ThgPu9hUZwcSjE4O7X5L2ThVdh7zqCmbBj1ZOsXEnknKFwQsWsIfI2kDE73eN8Bb
NC3IBNyaPZjjM40OUuCAdOXdM6sQtSEwyqXoMYHEMPw/0XsxbsdjiHh7p/Xhk/veXl7QGH46916q
DRAXWpTq/DcN+KaAxx4dxDzu5GYOzVlAAGd15mgFeOrvXA8QRpvwe1qJ5iXAW0PCYS4IEBJktOun
cUszGXR8fX93BS7vz1WEghHc2hF4tiwMU0ihDfe3LLuO79cL1fLbg7m48O+waoCtuBk4qLXCYkXD
ytk0eBSQyNpEccfdSrKhlCzjh2bXjP1F3AKl6kGuROej9RjDbE9iH6O1qxIQS7YEYNW1/XiEo2DM
IGQ0iRLZEF4WkXd99rW494GPxYgxjCWqj9L9LeA+clHKkORiHXm61AtIcDervuuLCPjenQ11jITC
HklGpr3P2ROok8/S6JVgVD3EK9NwpAG7RKJda+V0l7xSy4PPtV6xYgYGrWXLPdSbo980WhK064rI
HC9J/Dna9OBH9VeZFazs2LOndZ+dFDodvruZxrfL+I2skzdiVIKHehQQeqhb2ixQAIJC6cvT+FSu
NbCsnYhYc43cosbIPEP9Trd1A823F+tG+hvJJCvewpjte6xQ27EhENaIbiXmTcRVxu8OoxORO/lk
f0MS91YL8UoDf1bjY4VZQAiSJ9V/OB/IjrtW1kllb0KcgDO5A02laKoRZ8SPFBmRkdrV3p+Rupvp
lmvtdNubng7V+fApwapSBRHwrc5rFhJFFFLnh8Ca+po2cpeA6Vh5sUbucRdL5WR4Y/Q1rr16ByK3
MnkCr9bZw2DHvnUiU0bh2rhE79tb4Qj2kZCTQ+YVamC65NM5L93A4nE7HkzWX6HojVJB7Vcro0R8
RFH/jw0CCQtrOGTaDQkFOxzMMSfLBKyCPNLpMXM+V7BmWNaDKbBzmgsBMt5ZBRjGb6tdCPSdydOE
YKHJBHsRu64N1PQ278uGXoU2QzZikzjit0GaMOdcPV7FLHwhMOc5FbACRMOWqFM/ktv6dsJAuSuw
n0PYBXflo2osGZIC+1rYgXatE/dhkzZX9DoCJQrRskoSv7deQEWtVtTEVCCMEZVnS3vNQSXbnckV
WGKVYQ+OD4v7IKtPugQ+TW/BHKgbRRVxHfZa/OMLRM5we40dPTeEi60afbbzbWbZe0vMnUj1KxC2
iCeHpG0fFxLmkmb9vRzoxqpMK21uTE8akMY6Rlk1Gdu7YNQFWzryAcLkTpyG3hKroegBsryvF/kx
luPkBi01Yg/PB59vErOUKhS7GutOcN1je5A1gP3iYZYgsjYPU4JH42njHRgS+vuGXl9QdA9SEQoC
GQWy/dBwOGLx47HeuiWawVVQGhJaRFISdbYkmZF/wYr8rNrkLA5nRwGDKDZnfHeSxEqTulYh3/vI
zgxr2DMQxGAFoRQRHvb9jBT1X7vCD1kChjPP/7jBU2WVDAfrxLoOIFJNODkFZb5kxYOEOdcfK7z4
4FuiJQNL1gIUvrKdNrIbwh5j+NW4oDj+DQKqOpAQRwjxvdGb34FXpI8ooDKgFUT1fHftkoXOqOLE
51Y5xDYrx5T8IUkB9Me6Ynp9wzSgJiCWn7E3x3llH/833yRhTg5rcL11EuVFrZ80y8OvelsUB2Aa
u2HvieBHGwKxsXZMDWgcWreON5GmKjTNpVlX64ffhHwPXS/OinWKoqGqBj0ZW8Pb7F7hlIBxTJw3
6VcL9cqcxzrXp7rOS4vfuaqtGO7x4f3B8VT3OrRLvrILxvhQLWvmyaQhe8waR2F65+/I/UJYdwNq
4QoQy4wX/1efOL/Nvcby7s2pyCwutxfloNza7eNJlAeUvC92MrHJ33lWy9xuClfFMevj/Z9PL4Va
JZ9nPUQQu7TJ+5wf77woMxa39mr3bLSRQ2ugW67AvXE68YD6peG9fbGMm0ZvLUYXlhvjHbBAYmUg
xgKSjz70WvOKIa0gm/xsE5TNwhMdFoTqjWFj3LupftdJ5H91SJbJRLPy9vggDWvv5TPwn5ZTIUPC
yJys+DxFFksqEsoB63CzL9a8TUL9YZ2mefN/INzrS9uy1arMZTvWnpZT7HmzwjXwtVsOLp8vAtPQ
WlXqQbLHHyGYGVdkbxGgjX1BuuGsjQleZ69IMLlopax4k3WTmUBv+lEMu2Z5MwDFxucpY/sDa2yh
CljfrbOpXJLaLSZ7VIWQYginl2roVNvUHo/uIfOMuDoN9sfvfpneaoXZ9Vay7Yn5JCw5gWAxidY6
N9Ffqs335xL07+feqyQrKBJG0hbBn9SeR+oWHMED7FJ6sWfUS7y4rUlbQGERJHtp27VL6XLV9/RF
o+M8QIadD0WUyqqnpdiDPWD/3kMz62kuAe8g1xigCgLj6gla2iPGM8Wx8T36hxg0pJ7cXpMex6Ct
4HEzs6to9n8Wfr1gLa8QQoi8j8OH8PtDlFsIaL2vOQNfJdkgKfWMlteS7gEi+SowZvyGlJ/8hHMA
Rg7GnwseAypOH+kKySSWSIDTX/Q6NZrUFn73TBex7Jc/2vY3zj8MOA40wdTvQoCh+7a40HK/L53h
I3ERgVnxM1C5S+QukyJC5yCSV2PGySTMODK5ZD3o/DO5T+QIM4O15bED4JyoCxJRjgnuQaev9JZ3
PjB5yB19Itb4Je3DXb6tEz6IZr3X3vqfFJNn5WRVfrx5c2Isp/gZyTPu2qzNqNvjLbWdCF6WYp2O
kU2wZo1J9a62hYCQgnMOHbW1nY2qbM2f5DEBtlqI6pVXxlV8ydRNloSNbdxoObCJQ4mgttWcMkG7
my8NsM06uq+PRR90OO3UV+87lkyvH1r3M/wtBfb4odi6XnXz7JQc9GC/ZE6rmoVpPhCSeD4hKc5l
2k0IG9Ht1iaTFfpL7BwE+mmbEEwTeFEGUqElj5OOa/KZ4V2ZSgTrVWaS6yRwJE9TUHCcGFlvMCdt
+joC/fCVhiZLfVApWtWnPqjZvX5mfZMGhqAxF3JAcF5Lnz+tnozhhoYcLtlugBccIdjg17Kq3BG3
1IBl8lHNQiWc9HZxmIhlyMVnCUbBWXI4AMicaKgqc4b35192YBhIQuA0a4dhl9Wus0umk0Wjcvoo
fBIYcXVFxDPJOrOOTer20CteFrYuagZTlYHkmx/KPurzsLOgoxDKxjlbTzumFsqDV81gkpu5hiG0
DrwYzATGbCqgzXqR7J0n6/rtnVSvk1KoGcB3wz8dogS/VDPI3/M/WhjVD6ARBm5rp7M/rF9XSTeR
Z5zC0F0Kfv8IE6FVnwUUCz24y7pUOj5sPhebJ+SE5vgjWn338Rk9I1qNs1HpAfjtKUD3ooEY1TtO
gmTrg1BsbZB/bKJV1ac7IH8s/N60qvKuAcLW5wf+ruLCH36YCqAanlzfqbLUuzDbuJc/+TMs6OmD
fXTQE8Dpne69ogICMLk4hpV9LlRuSEO/z5ssuMWYJDMVUmwEVxRwUQ90/qfxRoTpCp2NEJy0Bb31
KpPwLhejxWvJ5BveGSo0uxspK8cbGwNm98PLV1hUeBH5Ic8fFmuA/7C7MqrBg8hU9DgbWJwQe0/7
A4GUGB8S6k30vQgE7bK1tT9GX8ftw/cbGpSte9S9WMrSz7KETuGkPZ75UrjEGW7IsbhocaQIt7ZW
j7qaPainlwAIUEFUPglGkXgY6Gq5V7PNbzP8azp/E1ZySYZvm03r70sKw/0pKFd+tTnXWzKKsx8T
lCDKiO0u8m9ufkIdKO1zbWIF+MaXNtV0P7yX/+vy9PJDamlqnYMFfjF9K+RL9r2nSO97T6q8kiDt
zUW5XI1FYaU++GpRXBAAyau9SxTrrPKAgzbVfSxlpVQ+55Hn/zpAdJT+Cjzo8SU7gBPwmcZiP054
Kqbibecsi1pSyeEztR2WBK4CLgBSVNnmpviPtqJmSxfK4AUQ8xZkkc9xlIO/z7F0qItwJNavT1p+
wKdiKM46s0mXutvVgvHWZSbJOPK1kXXLjyAqTJuO5ZDUwyf6oOjkm4bjWGqvZ8CZKoojOYlcAtxz
HmKuqfMKiCHqfauhuEI6lO8xjlJjR1jWVHv5pe1NOogtQGM+di4aoTFO5AnzvgtWAo478ug3d7AH
mkLtbPuFR4bIR6APpavZuGjCYKHzn3vWtmhfnJGkw4a67JKyML99dgB4qDghyYbJv367ei0RvJqt
o3QRZ6cLxpW7IUW5afwef41Y+Ji3IT/TlXivQ/uGntYwIMmDit6nOzuIY2EFK3fdNGsplwqQJ7Sw
JTALWEGpM7wUMR0zuHFZR69KS99UjOllC9mFVKcxD9oC7rQRgMDl32c1YlM9ovuEWDx5GsTrqlmM
uZMwHY25naWhJIxw24nClrDDwPNsvPnliVWq++wpwNAAFsBxMSM/A8zhjS6/LRxsHAI/57uGANgA
7zcGweZIcny8ZYlvqZr4f6f0XAjN25eR9g3vI1nTabi16SdlABMi5PJNXch512/8lk3Z/YFnRjIP
DTG/H/d6FhjMcYz5PXZedRNT8D4r1/1PnXsB+DfTm8SM9Nspzq+egRioTgcGyPP6jlifDFmLBY2V
15dPypRgZfC5pmNIujiy2dH2BB+NWOpwbU2YQs3cm6YH1X6Aovl4w7sBTd7veoOxa08m/SX4g4Et
BmrDQ77dQH/NiW1cKLb+NgyYcYBgLgzc1EMbZh3tdbXFti4YYHFW8VFcdImW4tkB5HaeAXBgZsnF
9ccu/E7zQQp6xvpBJnsGNxIDInQdgQpbpFupaps7DBGoR6YOFUBCg8yQFBwTkJpOs09AnPkS4Abc
Yc28IvgxoWvfyovFh2nBdQ2zcTPjgOIOTpGgkAwBCBMbP+AVEmMCxe4ynxl/UvAVMs3wtfOQf1u0
nwwUrTDsVK7gDXJTMiArcK0yqlxk6GaG44HFy65d0i0btnxPW8Tt1+KWZj/72Uf6Ba7wyQFDG3kh
xDmFyZLxQXPk8SHnCCAprgD2n3QeNwBYyU36zJJLdRr5iIDyZm50F94i7MOqAIlxUrrJ2Yy/5zyn
RVXigoUX8wnzz/49KR6WNKbVvW0WIaFPqA4LQb1HjOXQO+7iS4HNaOwDTxPnFj5mSAFsP2zqFAdJ
GCjZVYXO7X80gGiIGHomMWgT01EBWeTaC9a1xSUHRMNX4jiPIbNt2G+ESUKG6mRrBiYDem154UJD
lhqXqkDT/0HGjhKQgs/qUtLD/T4+B2ohFkV53YXqqlUq2GSPfke2/TW6ojVQaI8C5JfrUMkqsKrO
gJpQRnd3eYEUaT7Ii19aHqtCoCm8JHF+ukRdf6jw0zZj+GHjbC1j9ava3U9lTW2tUTxnPY+zjXm3
MdUu0PUzh67Hm7PnE/aKuf4yViVStJEy0QWClWEmRZIfpJOxvOM/cOtxLNHiEW57FJUcLqPLDUD7
kAFpzBJTBuQfx7R3A/PVpRMg5wDrkdg5RhzvvBh1Y4TFDiyKyabWOIGr787GhUXP7P8uv+S+0Qeg
2vG3SK9wo+14An6SJyQ8GErbNtvCuRlqPrFYww1WZukhKEwvL7l2fJ4tkfFFgu6Rkuuu3peTRy7+
jQJMYyfRmeJha1AvyipjnIBD9gxRI5bIfpt9sAGiPj6WbDiLlK4PLi+/KxL82mCp6tpW9t+5PG8x
5V6gDN6BLMTW5EUZsaV9cbeikoyZJm5jskaArGVJ7w5RsLGqkGqoBXkTYE6SGOZ2lB7L1ajryidm
yi/5jEfz/KMzDdnf4QDxBYFvpj7WJfpXSYLawtSNx4x01x/gQjzYS4K8j6+dA9uocgg4HaNFqcL1
TIxuJhQUnKarfSmEvVJUeHYAQMCLwaAK5vmPMuZinXqpPwSZEcpddfv6lA0OyBT+hKfuTQRIoI2m
JmaEnvqigiR0OceSHqv6QhruO6694sz+BeQRGieHQnuDJWCg/kpirYSYtNxzNaVyu7DRmZ7PbviR
3GkKYpqtWR47I2lVIcaRD03B4S2cAUh31VJCPoYnGZPRwyVgDTSFY3MzJpO1USHxSkVCP+TI166P
m5jFSe4POIolCcbR8tYOpVVuxAKurcunSXxO1jryf8hTrK1537ZdZXw+VtGEywusZQp5T9oCdtCA
ciqhqvhaqlYIgXjlO7PFMI+BOwjq/w4TBi3DrDkr0JkwBQsjFgmcY3io0SYmVwqC8JBHaabg2+Nz
lvwN66sTJ5gttCK/9mqO/awlvFRz/Q6fXTjdFosqoK3HjhyEh6kTO5HR5+9a4b/9BPEESdLI8S4E
MLnqeNsTwcdVVwxveuzTrW0TN8/WmZQvmNX2SCpsRw5nV4JWJbO2S79XfyYYgZDI2Z6WzQeQPge/
3x0IeFVlTvnUKAO7qv7d/dv3nCn5Dd9mMvLVOCekmXMKTwGXi1sAXpsyT5Ao2YxDdheAfzhuRk13
cbpS384ttCUnX8tUZzn3fHmVsXBpREAC7G0pongzYO1majvJ+gVK/zblz5zwAIxskZuh7CHpfLFi
a7D3eGM9jqcecOoSu4QY1glvt2L2wn5YIxhB0siaNeUQ4SmJgFPy4ifHT3Ql1YDKVhSvprjAlc2x
SWz2T4h7RJ+MWpE4I+HtevIIGPJdGDAqUZyYQXL7fTo4301MvVWQP9iToP3fBRKbV6S6QF/2Jfqv
P+KXbBkGut2LX8iK2lS4zmwqvOVlrJjzq/jLLh09SEw89UJkmKeSFOdWpNywU7ibxQDREcGCMfU+
JGiCel4y9YDnsiLic/fwLZWq5DP+dzcnCVTLDG5AVWywGtGQyGaYc/AiQnSIRkf12Jt2PtYdP+bI
u6g+8g2Zi69vVInjDDKwtINtW7HynSjPKDh7u7AhVa/CgXYVLB4Rw89OblMRx23ujM8e9hgYfGIC
eUaoVWQ8c5s1l9vcBhyjBZq++i7194R+S4gzVFO4k7br2QUoBb05hvp7ADztgo9ZsfVTzhtmT1+h
T2fmio/KwmERWTtPwixJHK43xc3WFSdqmWi5X1gH4IUHvqIzqO2rYKokh603Zb0AbG/GTvc0iJGA
6Hpw+WIETXABUVFFqDI6e4mY6t9OGNIPYutAJBtn767/iy7uKPKx3il/oBruz4keNOMHzNV4Ez0/
2yTu2kXpLhMsfQFCclOVGlC26IunxLtEe7a1swq0f58vFWcu5ZrwrJ92qy17e2BjYYHmlwOoSian
2OBqIOrA69nAu73ZUN0UPTxpZt0hdNbWYRHWp5WD387BoYt8LKGljrvhgbc1VvjIHipXWyQw9LOb
Xz6JOdz85bupGFuWL7fJx61iQWtSzX88tcWzlmMrOUwRwvZIG4f+NOtuxT6FBYeu5mPSpAdBgwWm
j5Fnw0E7RzsLTXQyH4FJR8oytrtyoFBvPDBNTO41UW7Q65DQH7r+1AQM68i2Oax8c0BdiDXKUlN+
9YEwdGX1ZK3XDAx3/gUAcqOBnjYKIwydQml5nh2h+EQULKIZ803RtgR8Su2NUa2XJsgivtwdHoOn
QlN7W9uk3CsvHcKKSKtFG7+wDnGiosmKNMpchNOWlztZZ84bHj6WZboVwFZnPCnE11sk29QAZ9Ql
MeApa0nXGCWHk+cYiwWCHyZczP3kDC5DI7vNBiIZPIYn8DR6XEbeJ859iddsRqmAeSx1K/i/z9I5
RC6ugBBkULsLUVJnTOGhjos7XBEvf+C32+2QlGoMb38y2TkVMBuC0uyPNIAkGlcNGGQX6i3LitUh
rOGoSTL+XQZ82uHJ4MSFsNnZZCPO574l6Vjo/4MXhuORAnk5iMBaBRYeZqbOLfpLqldtwkw9hXxb
tMKljmi4Mujt67ETXiRfzbWTx4d+SDE3JStYKHpbeQxekGDU+GibeWFvv3Pw08jWCdDZ4adtinz7
qKagx4CkQmhK2leU2gOU+/h6ntuBkUvEkR+Tc33AlnrQYZ5WKvbwBJUtxlmDWgT866sO2/+wcTWf
l8FZRF153JGlTaO7pMI5MbjF27dWUMe1xzNuksiDoeflsN67fiaDB2VjUJCtjHMrUy3Es7hpwfes
VPo0KC1i2CGCj7P4APu1jE8ncleFZ+TAtmvR+gmvqxnb3VxWQkH4mnEjja89z839q72Z4ojn2lEk
Ae1JJZa6lA5sJzPL43YzhCraz2llIGCGXStmXSWxs70kRNzQPLSNGPqhghcZo/nR3MwNyQYO/QeG
reK4zwUK++IGRXCd8QvZ9CJh7colubGt3ddMeFVG/QtWzfI8hATa+0H3mxYK43Z7y8omYASsa1Ar
F5LTfqN1hueeXjlScz7xCimC+4ux+347lZDW1Sd5mFg9y3K3nwd12/aKwTsUEYkS5KQQcYt5xtwr
+3f4l6lKGQlqXjARhn7Uncq91eW2SyeO73mSdxg3X0BnnXXFW0tlpMfEVDd2hKn2nRwOEHHPsM0H
L78gny1WzWvbzrVYmjlkpU7wxodozhutvcR4WHGA8D9T5FqdvWzTraD3Z5xJgmMuWcBBr5M09ktY
NG3LYgyAbhxA+FpYTHUUq8olqzvlz80vrdv9fk1OnDGgm79+rSJCjfADc5t0BeawBG4EqeOGlsan
yCWcyjFNkbIp0xKRnNRQOj3qDBh8cR0VeeCkJxR9wmjQrBo2pJjsbR4hiXY5uXFbb5OnpeTsn2i9
VHElm8MI6OkxvQIyCPn1dVP1x0ezXJkzy0zc6iXo3P/4TlUhaGEqPItgL0sWwOx3qcHAB0txStBz
MwFuVWj7B9pxdMaVBsOLgEXHqVKjbjdVyw9sTBYFwUBF2Djqfks+foGwq/1eyr6mDy0n9LiA1ZBt
lSHTlXmaOA0zKDEwad8RJ+cRAah5KiCZb05sX3UkhItYd2nHgTjDy+8JVO78HetooRcKyu59/nSY
TpXeMiHXXr2Satda678HUYFStT4GC7KyomgfOfwQJjln8XrcSywB1GrzZgiBS56/cJWhbf+X7XMj
bmubPMaQl7UHrXO39dJe2qvyC3UZ2SpF2eV7CezTaJpxrBrrOosvqX+6gOV+tjkxW1mcRrQb9fn9
AiGALSrSy8ZhWsV/OwF5N20QTgNxNue2gm1g7mYfkQJKmaifgJR/BU6QgG4yYxOhHGjzgOQSZwYq
P50auJep39wvRZ5YO4EkjBboJeG6s9LSpXOJegrznAOj6wElaC8liMbZXgMkNaMXQkfon/jhIoml
nWYQfecaNYfO/XNo0b4OeFRrQN9WLEKd2x7QNw9QT2sWp2hMkWxSKh1SybIe1rKdnmhrGDhs9qb6
a7NwTWAE12DtVPjC1sX3t2QeWIgoJ3iVsUTL+WJMNW+PVNvRxwlXNMMjlVRntfNWGRI/zMuG4sIg
KHLiVR88qfNPIdO1tdZxfuaZNpqDw0+rmg+2FmCC+Fb/XdjWNYWE8RlEYlYIOkMMmFJrGRUONgIp
Srmh9NRdgl5StuIXtj+iAL7h1CEl1eoIL8f0taarpSLAuOjzPX6ziw8bNyUKS8Fhoy+UVsql4Pg/
eLde7SY6r/56f8j0PHmeH2Ic5mrvhESIXBkbL50nmxITDs6lsLwRzTFMZiaZk4uRMopntTun4AS2
UdUEAgrDr+Hv+d8haSdyoX0fPClAfIYgqXH9Zf5dYUUBp+jUO2xi18kNVTZKZwfivjRtxcF9PfbH
IGqVMXAB2HM4j/M2PtxKH4OuvCkA7IVW8GuDfFmnvuM+8SVSLDXerXubjSwA4enrYPVMaZf9WYu4
u9riE7T2yIxS8MjisqClZQTW4s9Ey+vjFml07x2N5Riy+udmtzXQqs+Xp/MJbYfVAYR2PSdIVzdr
WB0wFOCr0A4m+GwqqslAYukwyYylqMTKshQUj32vu7FQlBan71L1JRYSsoPlVSLPuxOf0jIYVza/
aHGX4/Mcu2YaquoX683dzFo/2WwkDSkX692gr4eyydqXQQZxAGQX4oZy2VB63ykL4qvqN6R6WSwr
ludnQHCLYMoQ1qfeeLWl6cHTRiFKHpr0XGc8IquoNf+w+A9t2aA3rz/vaERtwBjfECGtIen3zVE2
Q6bHPYKt0qT7cZLclXYPVdLigdArtVZLRrRTwTJ/pGFgrrFhIU+nuIxq6qbUiMw0aOH39FLswCV2
B6xYDIdSNQi4/VY6ru2bGjPju0SRv4dms6wOPQx+LRX9qIwSrQGxfVEHxOLKNpQIH+TRwVmSl/HF
5lUeCeZid3OfVjHd/cqQnT0TGi6oPt4jVl4K+wMn2n02M8LCLBQHc0YDUrlq5cfj8lUejRFDlhim
gOwUkp0vSqTS67HvASAtcoIBq+jPgOWSFVeVS7yWO9/BAl3ydKwYFtndrVL2UzP3siSIz46miKET
waN88vEIer5c+pPtQuOOP8IzVI9tI3oKLaumfHPYlGseJlMBVFk9SQ/Z3ucQLpL54af6FWQrtIDq
BGWeQs7w56QNz++T2FBZ9O0oERbUDyQUPg0eHPIL7e2Iu+D33OsyFcR+ZvLdYo7TOmbMBcYB7geY
GAYoxXyrzDQ4M5M1ZwW2tCp78vtPi6tGqYvSQSNNeWIJoPsGyIrr3K5u/4ZL2ZEPlBG7zRUKXYff
DB5KCodJBMcx7OCW5GmrDRGMs72aaxUoXkNPsw08jQ/FwRkOa9vde5peJSosBprU1a7ZpqUVpaSh
ShKt3SQtMbiitxm6/2lX0Zcn+l2lQubiHqRGT9es3stPiFa6IlS6SI7J2R/h8OvjFzByCAld0pJ8
+b83ou7BYnch1CZUv99mrZlpZlYO5G4h8vI6cm2F5jpDQg0GXntrBjW/jjVeYx5mFzb7hUzb82MX
Cki23HUUQr6M2I9uNv+HjooIgUZhNbH06Y3BXTEGk44TbDzDmUsVv+lihCpEfEKLRNdXWvYsUCX1
bXBsJp7LdpVS0VGeRGrV+870FUBOulPUO5hHdgayU0Vd1pBn55monqAku85IQCcWIAuFu+/4aeGI
31KykFL0GZAiKUq7aczdo1W6W0viZV3e1A8RPIqJzVlX+dZ6q6oUOFQHjP9TrCnGJhGJ0wWAorhD
+aWJa1/Wz8HRCCSq+Bj00UyBqVpGxvxluH5NxkYzR4nFtgJ8UFgJsBPpaYbJbdssYcsrzeSshYmf
NvW9ZOwU6ID7mjRxo3AZxXFSr3q2pcKdXsY0kVBtc0hDsE1Nsm8Yu2kSvaXTDb6ztMQ78yhPA/Yy
LqJ+oW63HQv1a0pX7UbVeKkS+PKdxg7lKWgLkl1BkKep8Mo0oN1yWgciifXqJUdnH6wP3ayra2iU
xKZQzSySFS1423F0ZeKMbJrksqoODdgmYE/66Of81I/pfcjEufQLvizNJIIa8IsyMHxZd/8yUGb/
ZsnB/yNNPpqsmQHHjs/h9xGGUKecPPIoW6t+QQKzQCmdajOh+hs6mUGTHTKwZCcBfMImUZZ/i5/8
2coeDEPzI2RkP7dbrvoVRcHtFJI5XiQws0E/8ADgqMc+YanqQY12m5mM8zFPbxb6YFDMHh522m0H
3x+KD2Anusz8d2RZ9ONvBobH8HdOC76rZz6757QYa8zSkYTCvjHXCsBaGMF3VGcSb2hVF/ZYalNp
6hcOa56waHBMcCHHY7lJN2WlkPozEfNrofLoQ0zqWZ0ngjNoCtlX5xjta620tQ8lyABn5BgmapwO
mJpSSjFsPV5NKMp9bwZnKy68wW0MqIyTRf3265WRt+NVt0/MpRZs38mmOE62y5vYLpt8Okbho/ae
vY/xZ6/sKF8QjvTTFDVdkReKPhsGQ/OHyQ0orADKmxMqRDeY5z/TIPZGlCgsTo4wX4CDhsgKT+Wq
LzoV3TKUqBEbK6WsmLF113uujWIBWhBP3U32k13elV49OiayAkXxrGfEZS5iND9ijr4Rl00SFYRJ
/jkzSx3Trnxes79KPwvDOBrrSEv8jgEQBWcuMtykA+XlxK7bE0M7oz97H1AeXKyQV8Nc/ZKNTxH/
A0WTXlSmxmdCqTPlzE2uckXYnF0vf3MfB6cfNLsx1T4EsDP2nHMBuq/xZMyR7vfnzg8vsenaXLPk
2tJmoVpcgqwSoV7RSDplG39YRq1aFoWQvC3/2sNY1VNsKuOPJTSxwR1yOhts4urb/4NdcydWHKjX
HAlVo3rRkVfxeqk98n4QNE7Me6ZQTkRIVMdlrgcNaiwTdiNCkmzoxEu8J/e3eb/BC1/Uj8t7WLG/
a0sMorW8Gcievekxnx609a4ESM+/Ij5t555UnaFCqhh93RywnN9a52cm6ox/sd3Bxsh49k3RcKGU
XSTWNa9GXmuSpCWm4ZJ9y0XwruiImmRmpMyQZxLkuTOnKiZKUL8E2sk6AUZrTsdc6qfarHzyrbKM
84TvzsD7654rjU+B0AqpdYIpo4g9zxtrGkacp2ZqniC1uSLObGV2dRj+V9HcXKq3lC/CQfjgQJc6
2psZ/wwA89vZIez7t4Y2zqRCttTJjyMtoAqkFQKmQqUigdk29GNrakEybVfedQUuBmvpc8WAgauO
6qxD2CIOWDH3s9TXHtUOZvIuP9ApWmVivCHEXGTnPCZz8Ti35UKCpbqgk/8llrPmT+oZjDlDZrzQ
5qMzAn18vAutl6QsGD7tK0jrAywOLEuqOVr1PqN1Cgt02e46gpO0smNTwY4cyVkj9nnsI3R+EPs8
IE2s9PubT5ei+CIp37Qx297wDlv/rAptFkcmOlm8lD9toHmDe0pghaZEg78y1E0KXYvpTRojV99P
YAjnGmh/XNCLqBVQzSlAVQOMQDplcjJsKsBaAUQTEwuIBTAeMWWG4XwghHOq5F5KGwVX7UVqKbJX
cD91C4BPDz6c7Bwn5t+S6CLZWDN5y5f7r2i3ZmRx8WowPXieKkvtBT0XQRDebiqAMpnJr6PQblpx
IbeIwHncZd15f+5kEM685F1K/aBOtDlAS2JFuRQYFsRFAGevu73eJHAXfSdkRHTuT9nXrjysH/dT
wuSe+RRS4W+Ort1+MCwao+zsL0+V3Y5W5cQnbzoUaDnBz0HVBSKDAb00/ZECZ+TQgePEzTjCN+VL
BXLeD0yMY9hK86V7wNwX2S8B9A+6d3tJWplM9Xj3sGpBdXRlHIKGup08QldQvfd3IaYjP5haB4i7
CzmJqFyKKryFVHu2rCD8pplll/srj+H8kfdpfEBAzXiYMv/mKNLhU3CFymQzpXytCyzhmsGpHWxl
Ts/JcOAd3Ntk2nq7SI/83dY412lgKp6zpcAS0UOHZYlVzXJZxTxqGZuG8XaU9y1SIS5W1D5fRpK7
bg6pG/ms9HBs5gUSyYPUC6LriVFuO1lwxCRY7bO0WrB8505Ch5kow66U2UHpWzvZRmgrOwiFzPij
PWuzoaA0UlhxFftxgaGqVfzW9O45rFHq2aBt4OyH0/vmQ3E40IcnB4XG5YtiJQNQb4syYzDf/QSo
GxHhix9lxdXonqccwwKVQMjsiYxDVmg0t2o6ulNNJv14MDW38WjQRHR0rS4jBTIAZ4Z4IpmHmcy5
f8issZgBg+zZM1cVcS9LGhW0+30a5VCwmc1ERbfYBt8mcDMrRpDJ+oI3yNaMpQoJqWXhgkjNb+nK
L3ESp0yki0eIJY17g0tSfdJrPN/dENgYFtC92OJOLo2RQJ27UlArpGLiI62a4UmdmtFsCGlFndix
fx6tH4Q2u7GB/ig4v6FLy5Yj6YS8Rk8glZU2sle8MUO6uUaS5H5QKkJd9QioEBw50tAyM191LBMf
nrHY3LxX9NIrr476o6h+QB9doMWZNyDvOJxAVIj7U+8+X7zHm1s6KqodPqghG1Vh9NGDWc5brwRt
b3U7W2K2meN1CJcBCylpJcZDYcY9w9dnIjCQoRrl7W3MNDXSwo7J9DjcnruVB4BS8g7l3awVwoQk
Q2Ekn9di7+ixsH9p5e/zLEjzpSXrCbZI2YAfGO8OFPEiPo2oLUlDAgpSKeJ2G3+d51iJK4uqCkv8
DxvJmBFBUmfovyrkePUmVsc/RPMA31mOIhLLet+s5TedAa8TiFt2NDMj76nHsNGTJ97ojqhYSCut
cUdoWi1T21fZM88pgW4yL1DYXoGth5ePJa7VrxUOzI5NOLtbZlLLFT6Atp35kBl6X9+MNsCuqEjx
TZxyfs26w8qkaYX1W0+TgBFhOO0C2TG7+L+1GXNyEUDsXl7C0WhNqGcovb+1AFdw5Q1HEwjnlyjF
YREJ9lt3pOaP9pe+9wt+pJPYgX8XLiU7PLkyhiUbauKQxhKRkjImSI5M+jQ0YieuDurOd0u8jRpv
EyJvxbHmOflMXCTZXp4o+2q3ZoR+E5RfP6rsMiVI44IqFOlg5Ri32vYCkVSrf4gufX+cWc32kFWq
FvlkbWXdhUfa/noMdAKbD2+WQ7vB/mklXOD/d820DMObcpo93Mf+kx6B5bAsOnxzGY0SsSFv8tmn
8RZT4XYzgZr/q8YzpP7MPg6f6HePv51+faftt2NIFDnnTrLZxM81/bvOECRgSiC4Yx+bPVmLQ1FR
y/1FMfURlw+3PNmgKhdMsPQruB5A04hjL6+0C+A1meixPwSZSr5iL2o9FVgy5W38BNv0Gl2/cTTB
ynfwltLAYUl6ZsN9f92NeuGviqG4d9cDxKz5+Og2YaCWeLJVZRtM9CiQWURCCwbuO/wFVp/zNezH
wzRE1OUvWdlkGbT6XDwbE2iX8TJk4axiR51ut90xBg4glS1uNNRoKmG97ZdPSauSFUw0tCpPQx5M
iK0LEL5W2DrjnmusPI/o/56G3HWOBlsAKDwCq2TV+dUPRt6vSa2pnDT57U7h6J5ACDNVI9ZQIo5y
jFJCkVj2I98pEB6CXLhM06hgHtsHAJ4vwmb2q4w5pikdEqM3On3OAEv8ook4RtSJrynWSvlXuoPB
HktlAuu4OggiNMgB/glu93R+ByrBHFvXF/aejqDBXslKwYLyxoQtV/RycNu4tyVNLisYK6ekNCsF
3utSpIBhJqnjjX78ZbkedvWYtFgv3Wjyw/R2yIHY6FAlgAwLjQTbWEhdae/lYWahaeiCyPNuoUHN
j7JmBkdbA4m/8NZq9LrwNzraPGJGUcu5l3zp1FbHwV8qsJt2cqOk7mg8VTXuT/UlbgbWEt8Von0F
KjZI6ThL5Sii0mdr5VnGsrbCitfCeJwIRma9par9f/Y6VMikRkGsj50B73TBUOKcAKbOB6jK5AkI
tWT6i8rpzfuCmMN/dEpJvgJV7Tnjcyktool5olU1xwBTFKSrcVcu3inHacrWQ2GsbXZMS2LYMtng
xi1Axu3lG8uBB5lUZDaWoW3xsiuVweb5xBbcPsiqXbdfxC1ClBo/uylFETUN80VAeGNJrvK59+Vl
estx4Dp9kVMKbsQoj9PxoGw1SprxPpZktpoVgokDyEwWhdIw6q7A/KoeC9KNgCzNt5L5OGrmf2xq
iIiz9MYf/7y4yNxw62KLufHap55bOhLlEffSzOcbviqOkkT7NFdhQu+OXMqtCpk5ASg7Op8fikH9
t+aM74tLVM0U6O38CW6rufQKbUdTz8iC39lApehx+y1plWPOP8QgLmRcLOUFU2hNIUnueopWjpFK
QV9Q4XkDEEJGPzVBJUXw+jgrJzoOBE3ocKh8ez8TR5n6x0gCreYnZXUrWrTHP7xk/TIe5XCBXLL1
GP4aJU2wgLL65277fik8O+bv1SpDbgfR/KZcqn3zY8v/cUnSNpppml6KWVOhyTRl+nffAvA5lzdA
/RxbBDb2+MVC3WIELoyqb4hWSORCiBv3zt4s8+M6AMi2sgcrFTrtHS7r7CNkqhBLX2UmzR5ir4q0
ipFZ4cEyS3q4VUNMTGZcmOkVHuvqZXcmHXdoXw0dLX5zcHOQk679eBBsyVKC5j9KDB49KajjmebC
hR7rYnUBOtqXEBh/lraAhDAp2hh95ZOC0Gx2Jep0f2BJ7XTdxUMlY4RClXa4EwjVoszFtDBhsPXE
X6BW10c2ETVf/2tjDXjM7rGLaqYGVGqqr7Uw3IGtpegRUTJucOHboItpvoDAxV0wydWaSOArLLg7
BqwywSWEBNPkeombBhuCzG2kTn+TxsEV4zW1b5mgCZn4lGqe85Qgi1SVWSyjaDPWozIQCsaA8lYa
EKNCNAYp318SULSPOogwjOJD1otiGPOs49qEol7C9833wib7GwCMnkOM7n4Ytk3BBFjrAd15GMPB
Z3Mx7ioUJSAQZ0VIidKSsiHkYt+yBPt4fKAFaKZOz3cotHLqQVntoTW7zi5vCyG/Pp2yPlk8Da27
GdXsfNRblHmIzf6zNNChI0iILYAGKxyEnCM+lFRY6ZRKoi2dONu+D5Qr2Bwpkl1F2IIKRwpRvLSG
sltlZQRRSt+6j1GtTKY5eGD9LgwiHScCzyhczHlpgfu+sDHAWLrFknMuf/ajC6U8VmBgzETLQfBz
gjSbAqRLmEK4VbdIGzpVYUkWq82dOFVdj/t7RuKqIF45KMrlz/mz3YNoawH67kvGmunkPq7r7oGR
ySGgtQUE6ev7exOqjsO7pJW0zb9omH6Xt55px0HXM5x3KOe3jltOrF0v6UWhedjXcqaas2eGoEvj
8MXssnXeY+MzkAvLn0EkjthE9WBhP4WBGpBSMOY1ydqF4mjDixH2QveqP1r7r5FSNRoYmjjyjUUe
Ey9UiTi/w4q+o7JbKzwO1osKi3HsrsGQvrISAcGXLNiNbG43i7g6MGUCzXTUDUM9nurqHToO+8n7
47BQta9xUC2WXt2y+KJxgDJ/+MsLhfFmYxoeAHoOFK1wt3UhwNSzglqmD68bhbdq9CXY4UajTdoy
5xb9FArvPlXlU6KhcvHN/R+776a3GyS5KcZsDGkjPrrAcMJrp/Vl3Ef+zwCw8pNMbcqbw4GQp6NN
4OcOLSYkkk4o26dbwqB7Oqj2nZOISZqtpEadz4xRvOSDkYS3B66s4R8IF6aTI/uxcYXP1RW7X+j6
V5E5qIVZ70W+VnmSk+9Qqq0Hx/NvsWSd1ipeJXZyPjI0EkKNKq7IaO3pzX/T2sTDvanRHu4tTRLN
8Ykv5u9ZrsJGsLc9P2g5gxRMFlUeb8OQcuOJ6F9NV9kjAVlQrzhe7xAzvbQIZkbEqK0K4sO0ieFY
DAWVY25Kk1fKjT9K41yZBMjEUBhNBoHFJz5DoRWwGUGyaREMQKNK/RkIWecy4+NwIQ1dB1iKls56
umnLbR62u9r6xnntZR4yeAHumajUbJIzRg0c/Fgvz3AZfu/twEI6QJkW7/WZjZAJu9GF2h/lpsRh
L3E4vqWSJm50JelWwj2El53Dy7QBFS8tvcIaugqr4B4PggI+OhgJZmOAmtvMVxKe4ebZ9QviWnrn
GuKrWEfRmv9xN+uWNszuRTeWMejETJ1sJoCaiAFczwkWIp4fjslbqquCoWm3Vd3ZIyv/Gmh2Dl0r
IMjl8Og6SGh+A5UkWZk3ZV8onTGmVDKlKMIwfWynjjX5WRlIdztghyn/Vj3z1lQC/ihiLvQBBoLo
LQq4D2nldMOxvLVoIAlAO4LSCtbjEdN/8k/YzvHrMmHiPa2+kjknH9WfvqgF/WJ9GjXnMohkiBXn
1/Kz1TDTCA6KCspByqyM8cRhJAjaMmPJ2ov66zj/IoEB10pR1AKS7uVPjvJ1Mz46EJbx6MvE0QU0
ivf4z5Rgq1LuxkXtK4OWJ+A5rocY6M6/n6RCDWyk8Pt87nYbIrBjcuVeA/XPWjCZOGt+azOoUzVN
8uYMFDrrJsTP/oj9Jg9gN8C/wwA1JnxwZln7UOl56xDasTnh8k4ncd5sF2rAPcxNzQsZad8Tf1Ir
G7xF1FFIXAbtrZCjR13BjpodgYlSg+AB14lgQWCoMmlH8P+Bxbwf+Qb4jCnqVznY8FOSN/uudG7f
Ada+l4x+AXx/rOrKPpa8qjXyehqHbCCl2LqUMtgGEn4JaJFT72pnflPtTqmxw5VUJWXBVl80HZ0T
NuX+jn51MQuhgeQR6kxde4r+d/qL3XEvuYsujTVGISAt+UO09EgDCQvD3AbxlOJEU/JUNgCbREoQ
7WWjI6KjvvBSf4ZBIlT1eH1y+rkGHzxYVRSXek4pDqzvp2R7ALu5vdsf59BKA+10DveB0nmeRqBE
8Vr+ZUU1htlDFEWd7blhs81GlDAjOC+HURR7TMlQnRAERU4gIp2N1014FK/RcWB6HuDhZiRKyJ0K
YSRR8CqSP00U7jgGEEDDMMV95kqJ+jZBybI989r6tHiZGMX1zj8j6XSDZo7q4xJr45CXfaXDXl3w
kISwk7BJ6VzbfrslqtIHVRB5WtIsDyfZqE7Xyy3iXNJsF6yg3Sn2zNu2O0pQetYdjGEKECYqDj8b
qSbMwnHBF13Ko+sPdhF6Cl6aOd1yg7mm9TBq8BQGeZljIn96JGThQH8iGNWvWg62GgWHURJ+ML+9
qPTObrAvFGxtKixjQAMLkmarcPeWW7APyR92vYxOEJCXIaV+jLh9KfeqojVtOBlQlW2lFt1ORp6U
G+vLWoVwXBgqXrbIQvIutLGcDKTq7d+rpY0AFZgkOnSukE2gmBpesMSuEgd5Ur7UCwCVm2adBBGs
wzwF9Av1uOywA7Grnw6HRpNuKJnueggBGEgQnqs1Jx/QEpT8Sdw+8r+N8MSsOItQydKurfryLE/g
U2ntnchWHFpQ9lLWX2pWnczfIMwjx3yg/3Vf4Y3vPl3iJ7ItCnACVWqJ3WPU5YelbHe8Jx9TNIWx
bpqLy6YK95zOJQOkNAv7XCJhoCGN/xS5CfoVOqV1VR8th8r2b7v6sfOQStcConyvgdAPtvaPxdK6
VyWLjNxp+AAYGMjxhfDvZ2UIKJkfjDPkxUy3W40D11HI99t7sn04yXjcJ26yVtvNbguQmk/WfY3E
1nEcTdRp0mYfH3BZ2gQk7RRrfFemTps0L/ZK4nhC9/fElnmPWOJ/GM7Yct+0X7vy0AKLnjpgODMe
79JTA2nykqu7+0ifbl4SWkGVPqyEHsBg7HAyMQzOArq9V8U95lNA3N/0Ckid4hemMW20kqchrctY
D6A6z5XuKy2eBTSsllF5fTvHB1uZJjZImMhs6mBChKgupV2HlzU9dAYxjULmPU9iCyHpDZc26aGu
yjeyAdOcgMPWwAqmc4Bo/a1wfBUMtnKCIw4whhe/BOw53Gwc6XRrkFmN2+RAc5SoEexSMp6P9i9l
dQK3EBdNP9b2Unk6locCRjSBBS+YOJJjanVaYdBDMnSV4WlksHnNMrM9h8ZvXMZbJ3Jn0CAn5eus
9YCQo465k8b0nlbyC0HLqelyuoFJbN4goMfx3dUpRApoepKGABOnULwyRvReHqktypfQhPvnJr5t
obi1JPfOC33aTRAxGZZsyMEsHjhRV9tA+xInTbRFS9iacTO3ODNK7VI1300XlGZrb4RNyrg30KwC
sDMqjuoOJGfNr2fAVX2yDXv0YzMP6IBwMQIeYhmcIRi+H3PmxjNvN3mNgWY+759NYTr+J914vkS5
+vWHBYx7wHwSVnrcYJai0yZgidCyuA4eYWBnXPgpWwrGSXxPpezJH1ta3lZKTFnAFNu5Etrd6vm4
S8Me5UcVZ3SF4u1rWzrsTxNnslR3oDSaA1OrobXzA8QJaXs0Yl6ujuTK338vRaFaCZc1pk+8NuwK
aJmDuZJQ4o0Sw48VT1D5GREIw/Teeue3mXRbkcNpkazcpHf0BDsnxZoEVC9x9q7IeI108zkBozYb
vK/z3bE7wZVvQDmI8uCNcJE5XIMlXO/zRSvBITdcxc5W+qP4IxtYx5aFKrU5aThObU/fJMQMaFOJ
wU3uvRd4KNfNABY3VVnUp6tSKHtZZ7sgKr+AV6VdiMu/o6GJUfEks7Nu+6/Tlk8A8LCpJAENKvWp
F3YuQWPDnvhOlcku+gaW5Lux1cMoysf8PRAwCHmLInpseMS2pNphKWbd8w6duhcajRzj/P4UL2e/
eNyytmkfS5MekxzVpU0GIHqbW5cH49c2tEgfzT7m7lCb/FT+vsATmdBRi2Dz0eBT/ZyQexBYBk0F
W3pItWwB2ZKLn5mtCmtrse57GDZo23SNEYFRAZpBVhA9RrdUEsdsTjZ957ZcdPu/icPN5vE5PzPA
N+IRRQoU/GJlyLhtb4p7bjoBILdelZnZRHuVLeCtjUGs2gttt4X6zN575bSONrbYXdiqyzo/FTKz
ZeprTpRfuu9dIM9YSqVNKQqjlf721LdRQU5Wn0WlBDaJSV2rwA86LVMcDuM2DAqT1Wo8Qtx4VeKZ
cOlmN7AaUGMin6A6H7a1lS2pbPqiDrtgxOQGwWKtHgNFy4OXp6C5fBcckajFvIYRNuxfXomnHvbT
DUFkTwF3w8PAqTIrenGNxbGGvBiwMHvfdDWK8h05Zne0Jw9sldsuNq9JJVJpKEUZy9JQ5GTMzR41
jRnoDSPegXpgYopriqhp05ST1Rpq2V5pfFvLDdHa2zSd9rgqnjThY5+n0A2prIs+dz8v4JYnIuX3
NTzWLL3jjKEHCefgb6T2irtBXYQccR/cZdsfXbEoN/riNvZqjLqocboAO2c1VSYUw4QFoGiV6mVE
XRXNAmrbDbDP0D8mNIYVCuKIZNNsb9oojpgUxS5koVLodMZ0qIBuYk/ScWXYriLRYqJ8pylAt7nK
m47ZWlet2QomMQYvqY3b6g/rYbi1ed0xMYLidXvGSOGroZwfDDjrQQCD/oA4jQYWbyz0CIo1ENN/
O/tr6BMtF9TXQx2qfHJtcs8Kvyah3H88Bgg/8QTQCE4RTj01oM4rxqxIE6SZrpx8KCs29WBWAgoP
WpbyFut2mVVycITaytvEQ3L8/3Qz4I+hDUElxvb0H7Poi49uUE0XDAF31oCsAJVt7d86ZWdm5dNy
+45U9TmhokwCvp2VpwLgpmS+JW1Z/zB7HYRh4NTBi6aPOz1kIpCw5T88W3ke23GypRoOtDcm7kvU
hHMS8CwmiXTXD7lzOezSjPoip3zOkKZEqMC1bSpv2eKn4rsE/f/+SMAQZ5dLvxSlQaAP+Wa0RxnK
mH92E9gHaTb0Ahi62ksUY5lGH0/UK0QAkr6Pvi+hsmPLIZkVWKd9sIT5kaXOe6jyS7jH5zUJ42VX
lWOEZwLKhBFkeNzax8X8OaX6ON0towi/MgNXwco1kIc4B1KFyoFbXwGM2rgqr8TOKT7RqDsRIfao
zb0+HJYgb0dSUCWoGLt52n3MvWiP2K40HMjFjfyk0TrfBrz0rbZEGXCBqVlK2RjdPn601PP4kYfo
alwULx9oynVFPdg7X3I9HqFLyIhEm97zxKbPVOTDoe90Uqe7WEjIz5dImVKz7SeYIpRnvGpnmOpH
/PBC5j4uG7AWfsoVSiE16bQotmfNIxNAtsc1PrOMjYB7HTArIqhZrqShvCgtoXv4+nY8u4XHpfBz
I1x6Le769K3T9XXwPy0AyQ80c0OOf9PlXWSu3BLsLNPRltx8XSDvic9gHelrrDNxllH/gAVesf0R
8+Db4n+nZ4clWImreG4JY8tW0w+MvQu4HdhHFO6FETzbEKjHN8pdmfjjU9TNc2SdV7IDI2tyLdbk
KqIRvP6BzlAwq5P4pFi/MlRTx5w3KSnfmZlJjwWaCUdwhD5Kgmw1VI4xKAV9yt3GBYNgnmJJ/h/j
nvPzUnNRXg0ZuY4eIkoIpBzT+4tshHjhFY2CH9IyH93if/I52X758PNsCYfvGIyrqijeQyIu7Fbb
PKPta+GvMAB8hzCks9cCevfkgS8U3XV9xpbYNL43GbFGy+pBH1RKBAI1YYFUWplQHE96BC9iYRoM
22Qh0AU3YfQHQJShHO5UXuUwiTAvd6/vDRGtrJLGWBJe8sYbdCz2agji5bNfUgkbFJ5jAc4ewjDG
BA3ECupl03OHONx8p6FdJDLliGgw74lhnN3B0zSS4Nzok4iiCiIDGE/DAmnlsTwhrYWCAyBmiSos
hqSeMqxCBys5k6+w7GL0bju1tFkg9/NVgOTCSvvd/qs4vBG3njMNkRK/hPEDrSwz3RJdt59ItqV+
3YKFfLNEuQJf+aPwmAOM0HiuFvGfuoNNBF0P4N4PkxYjQLMuWuypVzdzHObXcwHbFtANVs0nNM4L
fZdvOZUQY5xvBDUE7Ka39rhodAaZl5LuUhi6XgBLyUKxat8CN5M8fkmhqQbcoMB2UFfbYKBwjjjN
6cTpPU9n5v+OvSmlt26VfFFW7DpExrdb9CpyWl8nYKvx96WysWDMOfPWDGKD5BeIOCSkwBZBfBH8
NoNKyN1o4MgybFFZg601A3xnPYfqSTezxridCkioN3NYKKjJk6y/5eUpUJHCZWY9YYN5DfKZjF4n
ikjoHDhhZ7KmnH6a+YZHhWaB7Tb1aopgz4T4WqEe7fEmGxit9PlrED3WiaavAGX2uxoX2Jyi/8Wr
jp9MX/TCkc7JIJux0Q9hcIGpwBwbUVt6Vgje2GJsn/+Qyx356cEhiVUvW1P8CsHmeZxxT7Sg7Irz
J4C+QT6+MT7MSMV2K2aKqN4CMiKQuqkU5kg201YmNWElhnCwhJ1sKBuf4vrIziObp3k94a34c0CB
c8b4MiusKBIAYC6t7j1A+A9/edOQGzuSZRvz8GrrLSOVwbWfQK5RVR57w/pB0S9xP47b5Qg9Uz51
GNqYSYitlZ5S3DojCWXGjziIeRpcJdCRJcKxWF5DCGb5WVBYCAN/KuqF7SNjBWhH5VLFJUCgrG2m
Z81BkWH3jcs0SmjGssixoUqD5FvQSjTT6bTyBj7eNMAylu0sqS5L2ZFKj8YVnzWh6l4EJXhQXPxI
NAW+kM7obrVqH9d92XQ+8++wDZAOvtDZlRyqtsDSjAaj5ApXQXoEfqLXA/2IdnHXYXARttGlqeV2
Nufd5kltsgs7NIv1TVqcWwCuoxqc0vMr06bjttKXIdol+XL78cUYmDSOsaFES6r9UbbTzLmK2Oix
Ukz4vw4/Z9VFT7cRbeywfUSnfS8uNj0YwQsMMksUa58LE4AWMpXFjrmt6iiKCKUjwL5vY32MQaRP
uzTaNiy9vHP/rDuS3sIp/eF72ft1fSvMhuEpQo/lxjxpQ4FVnB1q5bD9eDFuUL1VouwBB4X0RN2+
DaTwruL5bDJORpCaScF2groEqTOqjouc5wgg96KxkSH7fAp5ehg5uRIFMd+1cVvCqxPCeN3z1gsN
/4MNLvTb4fcLd5zWgrFYIIdgAdPC8AqV7t1Z47PE2asg5K3Mqj6NkEeW4oCJ6oy4z0i5cEreixaa
AnfIZL6hZSRlUIfkaqp2BKb0Y/pDdj7lbcQEcjtIfNHPLQK76UyQ3tVF/u6iVc3ZIVtHAafQScX5
5uua3R7yGnhjE/EOeae6WQQBHYOx55gwRcmuP3VF1L9Ypogwy/USeNfFRQ2Swc+dJUuMaaWHvDU8
qdYqNSkmcOY71SkP8PPRXfPbnFcKIdfP156FEJo3yWymR4/daENagd7X1KAebpjvUgaX2t9TsZRm
xjLPCNQukt8kZFsr+M9va4AAAQISA6k1Z7P/eJ/O+ZmsAaSYaeybWMZV50Owc1Mpp8amzoDi+6Pb
6bVgjwBzpT7EeFr9nWp6Iu++NyaZXNSCpT0ylAD9eZ12C62M8l6tvNsNGAaAzVuy6qH7eYzKMX49
lo2dW9vmnSDkw5lxCscCU9UGBlIMTA75SimrEDs3epi4I4NW+MHdrS5mShW0twoHdTr3hdmBFVKL
B4smrAFz273pJHFQiz6kKDXOg0/fCdmllmf5WLZuH1M0DBr3gNGrowyqSZ70vWiD7feLIoaC7jzw
Q44pF2lUNgkhr+tUWU72Q4NdFvh8DSup0++z1+J65RKe3bBvD9+8g7XYKlD5oirioJedoMdEbhgz
zt3MaKpEWMVcJBijnQNKPMp0WujYjN4QhDZatnch+mQqVV+zMHemuiShtV81Kt1dL4ANKttrqdfW
FOba5UWglOoPE1PsYOQsrfiycspMpixMzCnF7a3jEW+0TTVdcPXz6wEVkvJJWxmdjIYdrczOuotW
8JivS2MCY5pwgPStxAWwP+2Cf9ASIaoQlnUmahd14AygIrwetsJxAvjd1QLYXy7BCMlhUu8Li6yU
48CFnSlExxsekTyOv8rJh9XzSQyY0klzl2KDVdpfttQe07fSLbaZTuXrG9UIJPACio5N6t8x/+Fw
Ur5ACznh9HOvHO4lQukh1wbBy9+NW+dP2xHSJpP55VObWyxYlOrHI7NQFBNWqQCq0zZUhGVtW0J1
Q1vaPV0cVKgoMqhlUR+SvChig2jSik04R5CfQUIAqhXac64fonhrzsksoq+hp4vRpZ+dNNRp8rN0
xAzV5nGpmezXsZgl1BusGT19MrA8bxQiisWNlcijRbHB1wDgDf5bxDcZhLBLuHnnCH1NBpXskyVP
k+nSpcIE872FRrxNBqpr++7/Wg6I1WIX0tLRYCYnpBhH1OJlLiK0IRENnIURYdqDSpFOguIe3klU
+EkC8mVg6BVXqUGs/1bT+5uKjHDUvEHX0zCT3C7O7kGXxHj98xZXd/XPR3mjP8oRf3sUBM/oVawv
S25cz1aPOR5FCEW/AJ0q2mSMX4q1vrdRZaUG9nmFNZ4OPnVqHs8zY6I8goY959Eqr+W5IICwCxLY
zrwva4FYeL+P59tbujFCrn/Wh2OeYmGukyNVhpP6YMRHq/IPEdCSF+3V2i/aEvBCxNxQ/vpg6kLW
SnXO4eWVmZHMsrVwXyfWLMrlBkD8Jf2arMQBC99yYyEXu+updgAMK2UrMU0Ndd83YOubNjCxKI15
qMu0x93aLoypneG6vSph71sRFTsQ7S+BUU01PZ92qWXiW4qzsxegrsMeniB9kNNLimQ+uk+oLLDd
/EgDeH27i2ShCztHz9kQ5OmKNB3hUeiHuFnNTIHha5dsHv83mshNjPx04nNuBv8lY2qgoWpUZ4sq
hFZmHAZ+26wbfI/ABOYJqDkvfiUL1JPxkZQ3zUAgcHXFQFt7OUftgZ1PoEKBaYSx9m+CwNQqYjbG
lR32KsUZ6ldji2AvrqZbEkhkAZsA/JE/ZCQckzmK76H2GRnO5/x76AFRzjoZ0hEoaeACu8AmTjPR
/awB549BH2NfTJnmPgidJMPvYBADl7WQmi0RUbNftGkQC1/QN7XZ3hLzh8no8GRmSiW4Vmg7I+2f
vsvY1DQQqkJ9yqAziMk0NtqaWIjpxvwwDHXh3X63EOJFtPjrCvMy9EViJpsQ0HsNGyAdCZtEPt6F
WpOvSvSfjLBRuOy517EsNq7DLaeTCb8gBrdKuUZoY7YyE9Mc2uXIs2nddf0+DHtRLv5vs1UedtXY
VQxAHoP6bZTzH/5CNDW9QJNM7mBmSYgw2qyFP8hXmD3So4Z9Ax+dTl7VehhNJvIOybNTBYWHNpVt
kTIioCOJuJhd9nsbpMLrN9vplN+n7HSAYwR7zHuenp31AqTE1KrPMUrQ1g1oor/sUd6vFvwxOxAK
WyBWwFmnXvZWD4KJPKJB+rf+ZZ6tU7mQ3cpVMeO0VcQ+TYPH/UzNo8kwzDrj65+yx+1F6HQ1FIGf
L/qOEBsfDpBYLZeiodVbrX32Ujy6FUGwKTh57LI1Qmqf8yvaBPip2YwCf0hqROT5s31wyLL4DkZk
tQT5FFQu1Jqe35p7hp9yvjhV1lg4zdzvspAOf/QaUUG0OXzBlaq6rVyCa+bugmVAx52ff6llcxaz
0WTp3aDWSgz7AY5rqB3mL8O4hsIv1QhdtD1KYBtS4w5fTTutkJnlyoBAK1QsV0XoyY8BJzr9z2xM
uOXapGWxkQ8iFOUEF4CFw/9UMijuG+LVzlfK/L5uYXMDrYsE5WN1sWH2WNno+kr2yGB8NQap0e0G
tq739AJISD64RUZ6V/7oE/aD65jOlJW2XNTMPQnE1HCYA3Hm9nxlQfE2dG0po84FT/Tmlv8wniwB
uLqWhJKur7qc9mVLhQlW5dLpV9eWMywnO/CgwghE1rHMRs0etog/yU+eWkeyxsPy+6zYRgI/YSVz
C6z1j/Iw9Q8F5aoEUbY6dvRfItF3iXtGpF1re3Wc0Dvhbo+gLwO9Uavy1P4QwsC/LSKivpDn4PBU
tum9MQuDHGfLxmZ0a+0hOG2xr7WmIAYmuvQAPzqcOa10NA9IvebHEsv+FOS6f6TPohZ3u/VprIr2
cW2LKP7tkFZTVqtPG3RKqrm+5MDQdt/2XzvtD2eWU/+DqZxRR8qKuCQRkfc5YTQkAZ5JS6gHk4PB
3QFn9GQPH0QbQUxR9/NPh3xiFqbJLWibAnBKXJrSTSeEGLDoogscMfMpZDSZMC1/2rKF3TkwmztD
2Xa4lDKYlFBOzt98ajMcdZrsa1+LE8vwOll5J3b76aECJZzk8RuAuYb99EFTFkxM+VTIBrJXYrBe
oyJaSUHoQNhEoN2SztlcNlsXS4godyVGLcBo/u0NXvAsQcKRradiyMJvlpfRdUSrx874b2tsQ0Fk
YqUx+H2ztso6rDjPQY/tujxcVvXPRpYGnmleTnz/FRoIEXK8J7Uy63AoKe4FUrFPIQ+gtYxLB6s0
TVSspaIfGkTdCSlkKYQft69SMGInGAXCQm8JtV5xzqzUoyL5Cbrq1ivtUlkSvLSXr0EZuRG3eA/Y
gKYzPS5ETby73z3lUCbF5k2bOmPypSo1QEKNqgo2caf9g1Sg5VYSDF1vrFy42fcANvndL58KOJE9
U16eofHMs4Sap1dsbGnMTw7lgn2LNy2xgPBR+Hbef6HF5oubbHxVtHfPVHA0fzFAAEqsVJNE4IKT
uCnLo+/inogOmYlkE8VvhFhZc6Bxy83wFD+dXMP4Ac8MEI3QKTNMTJGpuZlcQRPk2iBxqAGVzUTl
Ms/Bz0RKG8zoa8H/tBK+yiDypsyUvfoWEPKBq+63fyy3GUWTG3YqH2Gy+MyHIOk94mzAk3VxhXRt
rnUmnnZmzwDfeEtkXxzM9YOLBm0b5R/WrycVJF7aG2OUV723Q8CF5KUmAl980WyFHBnmPEi8gEdf
QRbxny5y/2N5kzNG6sPyVWCW7lzHXtuuVYOlPNbDqaa47na/Wq0XvZUXCTbZ9X6d5kH/h+0RLqKd
3Tdg/gZJjP7mUxS/L4FfHwYvNxJbb0UPeV7E/UM7CpZ3pX9e8LV+yhCI7MjNH4Yu9+n/AE3ICKz5
W1nANPQQ00JLF59dSP9vjjXtyw9Ui/h6OHUB0Oaviu8N2guDUPvfAUWdRwWYabPA9AY9qtkyF3cT
NLV5wrWDY+9t1Y1rOfln6qc9bRAX0AGkoy+83iXrtkqDNwme4lq0uJGUNmlEZH2COL9SzQqVOhuB
GpW+i8MKO0b2CV/zYMoHt9iCrjhqGZHWw9PpvuCTRlvHi4UYTPQmiBHx37rvmwh0irTCbNe38roY
bQkloeJ9HamBDwo4ObqJoFpuE6o+HID7vdP3DJgX9KB4jOEfwB1sDCgwwOymbOe6yi9Ggtkmd+gC
sI6O3G3T7fL/1N2Y2lQeKp0xM79ubp0p+KEiPEFwRUgsJACXwBQa8tO6OrtGXtFf1AcIqemQCv2X
a9lLdnWrnvsa4CI6ifUNrOZJ32Ev+nSbEtCTLiL07FQxe3mJRw6oeYA2dtyws4h+KM6sSqMyxu3g
iKtTUBUHxnoAvt84BTdyQBRkmd89kjvisY1b5Ypp9+qjf2qGTf5Lqi/1y9kbZrSJ44tAu/NDDM11
NgvpSfzKx4L8pBHobZ6Y2F8iq72rp76k6ldRp/NhgfS8TCXviXMRB1fG6X3lJB13Yb8gXtRbYoLR
6oMQ5suiBWuFPxro9WKPZGm+2SWdGV/lE0M9geQbM+h6F8uWuZEBeCezvllaL8HeKeLEEa+IPyA3
v3E3lswckCljA8cFd0p8cmRBZIEX1Dj0mOsQk9DXqL3EKLieOt/vUa0xYHSi7HB/KiLdAy69l7fu
5LFwRCorgiKra086uxNtnmKI1Pu3G3Wk6WEcxgqqHWrUnjzKyy332+eQcVVoP9PH8xHNe6ijwuhw
3zUZvZaAWlZY3llAjN70euVF/cnF6O4iNOrPBvT9qyVeEPe02mr6KdRgZqskpgUJQvnt7HbE9tVw
ByIKrYfCmLRy97r2bpA5YSp0OgnTTgx06wIoxbksUMUtEx17FRXJjb8unfxwwuj5U4UCkKhDN79S
mSEAVwzi11S8AQtzXOP3LQ250MarSQCmGfO7xGRNWTB3gNg4Bs+aq5htHrGcLM/YPw10iV/vF7qW
RBsGf+cuYxzbbwkokTaYpQCbyEm7rNei+Ut/vh2p3N59vqMazI0GBHZcuuDYGmLxQjR108/apJb+
xEeXbT2ff0SENhRRvWhIgbRItF0GnRC0dJIlOEk0u2M8yRiWnODOTm5PShR6mYubQKPSloa/SvoF
fo214c/Xc+3OTX3deIUjwtJN3dPZ8HNPBSP88Fsqs0HhYKxOll3rP0FjwV32E76UzpRa8mxVZqt+
E3hmTLvVl+Wjb3ybGRvOmSf0I31Y20Ff4dHVbhCs14vfugE80iy/ZuGKl6llmXPGiGXas5neD/cN
Ye6t9jiP8EJ1l5jceyIYFwL5qBfCdhx7ZXWdiE/W9jbkFqZuPu0DCuPudzF4nR5Hg7SedRPygUYm
4DruBN6y08IJ6IDnlt2oom44dDeh8o/uTrJpgDhPsQHYSgwglLLlcBwHe+c0RvVln63flfriC856
Qepv7xzxnBK7iTBGd67LkbyFmCwuSNYVEw4Y4DPjpZRAoStRsrTT/jVconci7Nwf0wDC9UA+QZAw
YeVjH0NXxOE9rdfx+X4yKzWiIWyJCD14szXLZghIvwg2tEIk5XdbwrKxBIAcyfAt1ToG5q2BZ/Ov
5ZdGZt5nJmWdJhJAFhIlt/OZqnB9MEhkdyFLxnm2BlQTguMIH0hNgOla+U9MKD8oZxiWrEWnTswb
dMKIP4C4BKkpWF4sgN56u/WwNMVXSBmsHuu1Mx995KylX/PnWgNFDSUOU86dGvZmXWlXg3oLE1/D
v4ziE8YqYRGNmXBOto8rxKIDcDpw9Q9qON6p5eCHVPQxAaKxbJbhOtm4rhig9ink7Gh4luvaIw1d
MmrkHb2oJorrIzKw8W407N6I/JzEXwmXLq03iajff71lgRJl7bir8FDErDGYPuHyDG6ECe9xYmsY
yq60HD1MHkx3TBoB2Gp6aqLudy9wCPaHqVI2u793Isz+nAO+wf7FZWktDNPiHQNvmiWVDYpPT7rM
+fgysrdrMgBkEnvi9Jz/4GDzr5HrQ9fiDmwfcKA4RNh2ZCZbFcMwrM/c2hivmhLTW8OZB/QE19IY
4mcXL8Sahnb7qgpajvNti15k58rMdc3nZ7fohpvrNtCeGBhp26gB2de35gw6aGMcvpdtNQ8qdTYc
dh1ncYs8cpgeX/sfPyKs05j7PpWaqpwnC00AWpsE3FG7qvcDId2LV300bYROTaXC1unl4/cnMGTK
EX/AFa5h8IXaN1BE0GqdWZl6IENq0dmtg5xHZ/zQy5UEG43yGIPTo1RtfnQtEfCNIG6s/qqxniaR
Y/33L32YrCyqKgR8F7bxBiWmF3V56OgEE+GxEgPfe8Q9StrIrk6incjsfqctTTPC/m8DT2ssbJzc
XqT4WBuB+8RKZNnbgaoHwnH/oEvZ6MVKYiv63hos/hSbt58HF1raElgcRSu7/VwALuN6UuUi20e7
DKBPPIx/lT3T3QL1zGgf6QDgBgPaZ3R5DX2rIsuKlJfLrAjYj4Qmh0wsT1sQaiNzNz1mrWSTziky
fYdIy+pc4tz8mgqPieq6jgN3VaXKGn+c5UOeAiBZCS/hCGalLleojNe4b307h9iaf04O4u/0SVQe
zFYsI/v8Tb1z02TWY32sBkLIex88a2dGTAeMfYvUgwyroZkZDv3d7V0rbmEvM4RxYUGuCTptFXHd
0JChVsU6S5rFdMYIMsPRfi3AI0U6S1reeV08Ro1VLKScq0Pg6LqhsXtT2zaN6xuKJfaBdVvuCOyy
fLRH9sLbPf4MIMyRZUeXmAmz2tdLZhbdgoyfGt7gT8C+a8Z/2/GaUfeAIIp0Uhe8HKod0kFLqb3e
E08uhQRiwumSvcktmuvFSRalpvFPEndm54/8xDK3rHFvV1MrEBKSQbYK7PPymZyBdLmPJQoYjQSJ
bGRi9MDvAHEX3y81jgUV9x/xIelwlnR/r3soL18t5ZGB4RCBxk7T/IcheFSMRD0e9GJ9BGia/tS2
Vu+6reXYXQggDIjOQDOQCbbbY+pN2Mc26DKXfoBeIARv0FVkaqG0+u1PAddcq6zWPZuCULz5pl6T
QNR/3Rpu5BJF7/kIHEa6lA/2aHlCLpnm9x6a6QomO3e7eqHL02jOWoG5uVXR4Wq3PPoEkR+LNaTN
HY/TS5aLnTHT5F6S4MpWlsCl8D7FqgR+mDqJEEsKgn/R0bkcqaLdRwkqxnN707EPFsXfBQDDwXGm
iExH5K3OUbEFAYqU3rsi+lSaRm5nLOiwmfg1myNWtZ22LAQp8OHOvLswGS/5SmOuESfle1oP+P60
Dr1bB9oCGI9wVjHs1q12R+6ArjIQWq40TYrEOIvPiB+MT4UeZdWGry9UjrQHXxX0k58WRJ0jaDcL
+cNafRmxIDYYTQlPhJvFpzKgPabQ/yq8zVvUFvWOitbL1KIEcGYYoMobBGSSAXSTbWGpesLZYAlH
IlYsXnx/4UXNlINgFuNeZCRH7v3RCpqJkFVuV2NY8qEHz469QpglkhoDPMSkD/5F5jdNCrrGy+DA
HU9SB8vCkTLkdH4CTo0X+tjgGopUKwYZ8h7H1/TGdCJob/rITo7IJknb+6R6CEZxcHOFdutarxUw
Wh4QUI6gQDUirSg6ao7IlA5UnA1CYtFbQgovAWEhHbrpf1ntE0zcNWg5JFYnMrizXQ1yDWNppskk
pNMNP6rK3MmK7KTbMueKbF2P28JW3vq/x53dTMppGBpZKfU/zhkKNUw/+SX2L97z5+/dQMw+5o18
N8KSLx8+eHXX6JaA7LYOHyA/wnF4mKCR7Lti6XA2Zm1bM6LmhIc53F5JiC3WR+gFZYzqWnZfFU95
TIJJQArLl6Q6uflLpdxdKDWl+K7755hTKgciw+Dzsy66Fk9aC2E4ktYul6CCiZdbefXPMw/YVImq
6voMIHecwHPitG60LjzN07KdNPnkr+ss4AOdrtEbMM+9p59TEpKNFEBPHd4UWe1aApcqp0uA1xPX
5niCjATFMVY655nukBXErNpAezcf7K/4NnDWUHX2BEuv1sEuwi/eYituH2AG5TzVwJaRQfDquX9/
NhB8Wk2Le3O/dBICgPafZ6yyirIl1BDspCctXRRuTTDa/jUcJ9fJYcccg1fo9FyLGYJ7yprOz+Ls
4JTJoSn0zyYiMkrXd+xgXchqOmZvwPayvuqP/FGhGVoToKRFB4p9lj1Ml30uGF2jqDqTdy61o1pO
z4lhKOSMYE+fGR+URhIaPCtb9f3OZRY6qTdnD8QvnoKm2Pg8nnVUfISXpQaQS4uCCrgGElbzspWD
sbOFPMKTAZma/p+Uth3j3fwdTMimXUbrr8F9qAzqB1gKuuYj1/abDVtfd9h3c9qHMPUq/Vm4A+/N
mrqvG53Qt8saF6istGvdMCIjq8C/RenCoVH+WnbX2HNn6U6c0NAiQMDgMbM7WXkQVrMMZsuE1Nck
2YBYV07kLVCXYiDm5MXOUL8RZW2k3UVgFbPMazQbzTlnvn5ST8JVWA1dpTN/pRD8F2+5SZqWN1bW
sA67fBt8FDeA8Qs1plY1bhHqSMIybTBJ73ki1VO7yNFDwjcHNeLOSmUdx2/9yr1huiBDGrksnI1b
OamCZdzRYu4TBW+n1wA7XbkwlPR1v6P6tbAzRKFccKz+zAFcgHfJ2FUrenCgxVhWNe0h88foXmaK
NO37xuSyKTuWpbhxsnHDvSYDP5MizgCRONoZS2KR752ufABx3hn9rjN/KNijoJ0DN35S7InVhYjD
H/2wkV/+X/a3kOlOMJXpvKB4Z0XqmcUTrC371wuMdM2eNbp4pHR2uN5kpz4ZU0lbgLf8L9VQYnCf
9lXbceKnc1axOLG9HsJzMVrPJ+yT7KvG5THwBlH0h/woFbNDDgdzPkPSZbLM7PkgTm1SUMqYxobH
XLQf2yyXAU8UlG4wPzf+hqbBkbipK5+HRqn3Gwp7vubhdzkPXt1jTRrFnsEJpjRHsCpBq2fX7rZT
CbZtWQLGTr1B5kkgAEUcByff/DSxTzFQ+uF22A2teOEFHQAbEHiO76VH+FWlrFWW4NFeFVwWlHbL
fdctS/8wcEdK60Od2fkcZaSYqALCWcHa9167mNyr1WV7bXd2QaHF996EFU50nJyxiZOIaxUlbryh
P19Kdt8R5F0pdxMiW19+5JlHhm5ywoptw5JZpnTZ2DsfaVWV6r7JdxGhWcSKw/eFv8d9GNJ+YS/l
lIXx6mYs8EWq4cgm3OJIMQtzoOEX/+3tKYhagWQn2813sOHTwVT3rfkR0zWfXRxNy9T2KDKRDMYd
vpPWgfmIe48vtbfXiyORIBfwmcNvpCZCWZJx5ktZMV65B78A7DBLgmKn5iS86PpwTlQ5SI/Lc0q0
sjrtHrwjHRMYyvgN/GhozUVmRKul01xnBJ945f5wwtMO7o48Uje9EDzkoxOO7hjdCRYblJcUmMLF
UkH3VqBAyFoCdMKYjg6nO3kV14bkblkodrvsI/cA/SBP+UeMdj1v83FBA5EC4eioLhGicL/FBbBD
e4kRW53fW0ilEYCVYICJZfG8gi1VwvtadyqdhVlqYS8BZP7oDRG7vkyDtEcjNenrgHRlOYmtDySz
wEL1R7k6VSZk04TSbDlHDzprjJCj1hE9nL7fQKGl7/7mXILWdWur9J6X8B5Ft3bYY5YcDES0/xZR
zzb5UNwsUNlnzLGIrLZYkX8oKuCCfxLI6PBVgye29e6YC/ZoN7hP+9M/x/CAwnveaLN9JpRrvxLU
V0BN29O7QKfaMxSX0vRB5QPyZnr58qfYexrcid53+yZZIsHiQndqpymtotCTn4wPXN4IDWi8D+1X
6SDcCQIb6LFrEVyWUv9MIYx/+d1oy+rJC2ye0h1VKLFCSCe1YwtRisQ4O5KeMDDI+TP7Wbcr5x3/
g3aIkBBjBoedyW1yDvATiqb2fUfbFPdkbgRG8p43sE1unATGM65xuDiPw4/ktCoAisF3m+1T9IlU
RGcvAshr1On343VrfGktwI24uq4H1ecfZCjoaZ1eFboQWQUPjadKsZ9vWfXRWkZ8xK7GU2i0fCAa
zXlhOW132/urI/yyGuIHElytmB8TnBE897+yl4K421TXvbUn4JtzwWvBZg0p2dddb2lseBtBnths
SEvmf3xzAJc3dsOsEoNHFf7CuIsjVAj/osbsinIXvmo4egoVBopWeWruDlm5IJqPgkn1jEcj41v3
GxV76UdzTW0HpZo7cBcRkVNfdjI9BE5bY17Vgb1uWmOPDdCVd9OM7qbweNpQxpVHi8GBvRVUvFyo
fSOAGUY87rPnZqbYMR9i20s9z0EGhz2/mKHdtTuniQkBEMUHd7FOlvlHOUPHVjG/EM79YIRF/dn+
A1f970NnEEquTJUEaw638vMmwCu9ijS6XbcjvtOCfAL8MpAUOd2SWoa0qtw01kVoeX9gtSkK4clj
+wJLAXGFA4xKMKlKlotPAfJbukyZcEjcjdsy1rPdD+56MiLHRmVHOcjhtbHiPWywLZ0aAplkvp5r
vcQvC1AR4OQ9E4iinBbvbhOG9YQt7P1U8HrTLnqp5stD15pVSTmU+FaijbGt4My4NNKSp5vdX5qM
fDvUoN74wNsUt0lSpqfmpWhiaSuJ/D3BQRX0W1TudGP+g4/Qii25ePTWFQupXlfswBJDdDGc6v0x
6oiPYu93EG31IXRBa0P82UIz7tg8VhrzSLQ4BR+9pHpYO7GI1ybLQrmVDtb2FuJwYSZ5TWz3HoAw
YhiK6Xr5+G8CBtCzERNGqtkWRLhLy3/fng4tCiSb3gQXwKK/489QFo3xDyrqnTyHI91Ejg4CTY7r
fUl53FoPPkCf+cmr/wYM0CsFpLlIBzirOaeKXbUZnhG875V0TnA6zQZ+rI+JADhY7atSqxYUS8Ma
QsZpbhnZU1DFc4yt+ZpxARA5cv9Zxl6QKgyPVEseIwcnuto+E+XXszI3J2hoxO57GCTDQp7fSQec
X6EEy6N//F/WC9ftzxMT/2FRP8TN2KIzW4cTLr1xdbKTPreSRJ6kDuzTsIbtvi4g1j4I/XXSzMB7
kv7wGfT0oeMKNR5Fppja3XyF2XW26hb0WwTIvrTgr94nbE4c6u0jRkro7j+6sGbQFvzfORj/H5tp
SHqus1YbMzOc/SEuk01tAdbhFawgjYhVOV/rs3cnmYajgl9v1AgQ5oityIaX7BQJQIDAY5OhrXjy
94B8YziTKvoYXdxtFey+zZ5z+hXyWsvlLMlXihxo7XsVxQbGmsbpLogkRNOCLhjecfyQKH5wwjQa
41BS99i1ylmd55DMnyjcUUMdh8OjAzRK8hJ4ySLT6alubnEpu5lf3/V1TATnacR4AlgnNzka9x/+
f1mw8DSGRSsw+qbkHCWnpGfl6tQlOejIDl+bvBffsjc4N386xiy3szudPJLpNSw08iThAYi9GGun
Hxfyn3u+TC08dxp0eAS4bAN2GEeWxvWINKpx/l02lLeCN6h8MV1x9hoyfJAByPdj7RVSTgcHaV5A
EElVr5TJ2d4ZEje6KF6XJsagpzxCkyGbqmigHjLnr80r7EnBNwBUVb5ekQIyIP2qpXX6hLlZas7k
F7AChwuAt0e87dt14PgrfDUG+YQFj6up96ehi8BfGCG1tSYlUZCo7VmSQQHPfj1Plm/d0VT3wi0G
HCUjcFED6QqxaQqjlwVhukrPOX+i2BpyZSkiGmyfbu1hXREyRp4Cfw0XftRaBXRTaXdkbdPsn8OD
PidCMi3vSKlX4TmDnToRrT4T28X2oamCxidp/lC/lFHbuluy4ik4h7wc1x4nC5r1vbnuIYg2gKIX
kyXSLQRpE87Oi4HsSr+gO2YpsSWX7u7dDVYQSeLacqYx8m7bcBa9qy46rOHvQeqEv+Lg8ViDOE0X
dt6fSdgNHWJj4raNh7u1fkPPMb09Zgi0779A0hUX0jcvL8PJVlwtGtkgXfQMvtTp+1twBoNROPUw
B0b0YRno4up5TLZVQTbPoXN5ITUwr9xuyNgNBwUBFqjr67BzD91UFpfER/5y5rCaKxGwGsbP5bfC
JQjnLX8qlAKlJyCvH6pc5wfO3gfqQwycbHABFn0/RiQ0vDeNEWpnrWtuA1L6FuPtOJt11kYOLqEV
1jnTD8zudA7ORC3Pth1rN2y+OZ6lo/5Z7a1nRyAs2G2FJtZPcg0KhkyZkIKo+MMnja/P8z2fT6Sq
tcMsetScubqykxpGhmlWjDIqOFO26wH44hvh33xuqr9zpbjkblVVt8l10LKm1+iYzYineVkNMNmh
eg67P81Q8s4u4DQIEHodzHOuZkTXm/S2qh7BiKSIh8+0anhOt7JiJosL4RY+0BZ9IxDhqaXxH29D
NY9N+tbzh2ecrGQKid/qZ6fUXG0ZC+joHtiDcMc45zuw8zuIHgx/uFBTxoHLJPo2UbyCmYD9zV3/
0DuVCtSlNJj+aqC/GsGRv4GiAR+AY6usOchUPYqNBjq5s8jIng/H3P6+DoFjti/g7/jjTcBExuuW
7UHFSq2kmt+iChPL+NXJTYz2LzlQxXCLnra7DmGYA75eBmYQbzAHBE1TQVtWfT2aasRMSlUIiMmU
CO3aR8ahjfcxk9qPfi8kDnXjWD1eXvldUIbCXvvCYie8C+XL/vmP8tg9VHR13P3latkCxNDb2mza
CjJ9TRJuWhTlJD4bkDhI+GunfN6UpeUeScDrMQI9pbqjBno5ClaXYZ1sjvzmOcLQ9V1YUkUTPCu9
q7gfw8dj+kz0YeMQNRA16blZQc7GWacXBSnxc7ieYGuiZQ4yM+s5Hnz5ab9cOkt7MtZQUSikZxBw
dwWwdBT7ImuEV116dayTxtyKzSpPThftcEwqUaJPFqWk8LT6Pl3aeN0WFsknZEwafPzwHZF5k1i4
VbszHdC7cMkAh5SHeuJrFNshMcCmg5Qo1Ujh+8rO04jnsYcwJ6RDsKIFOlZ9VaQYgx1v0THxUb0K
iH0BRhYHS2T74EAYgB+fIJzI2b5Ex+DuouFZMLvDC+VYrReDeUsAFpq8l2M9SVF8flWZ3hLlewws
GI56KH6q2ecTrIM8k4Z+Vfq0vWj/0Sq4X2CitzqTzx4W2WT1lM7i2v+LWawWBbc+HXSkoRkVhF8E
GfCz5t44pNDIFSkSGiK32Fiv7v0RaxOMQo1NjMfQca9s2SCfRDJkzvvgl1ci4e+1k0JRYblmMX8J
pb/L8PdL7qF2EpUHrQnRAf58uV9oD//rROK5nUzKRyb6jcxYi3OwjO+AMtVBSoLSUbDPgRT7rdym
63YBmZH0FzNOQQbSeYVtVccxX0b6Y/nvFz0R8/BBFZwiIQGn+O5Cou8VOc8CedvErsnhxlFQ5TYX
LgzoJT19DDxMZhcsJVYgjh3e2zHxLyVf+oGNXYWAVuicdXdJJhb0e4PT/FFJJ04R+/mZFacQR1RA
jOA6ZdUdEoe2JpehhkvXfPnsdX4VDG+0E/BUsKIkPrBr9XmGpOOtWbHlgASvlD6AE5njGgVyUHu7
wbZf4p5pYMC4LYNPxc0gqoqQca9kHvrfFuIHzsVIE0S5/i+HANuJFIDF2x3oMNolJkTemENDt7lo
xRgFMAQxt1kYRK/SV7mQQ27XL3KjCV9mYn9crk5llYbGn+4pMJFBly7PfGSjE72WLTjmij//hOBx
8/7QbjJnJ2U6XRLSaKh30QPGO12KhpCK3wopiu2GRISGhY8Xrf7D32Dqdq+oPf1Bk9+6R0vRCar+
0MChsGeCidCuK/LDgcQ/hhAaKB7b0+FL5fKC4zcokSOv8f24nuZRe9DHi3sVR0q0Q9Ymn508tN8y
ndAbZ80hYUhrmRolqrvgtioMMTp5dign9mSt5RiI1QhdMgfgLh+4Urxh/ZUgY3tmDtKC4tcmhOvC
Vnyzd3ur53cTMpCdJE3dFc9xRN7jF99YMjdCZdOt7e9iLR/aBa7+Wa+IY72QMADdHqzkK/QLy6MH
EuWAYQ4R6XfydhEwUdhV43Aidbx1gJZIkl4/Z1lbXOqUP4Nj0ZKCcGVPF+mQx7AF7VOByb1EmWHd
fBWR/ppkH5RRtF8x0Q1AZ4eELVRaUsBPUhfE4u2VjLEEo6vznnloaiIq/mgz/UMpJKoJcylRs4D0
63gqh6q+4WISEoI6Am/9Q4HY3bURQDntBVYUWGCm7XlwXsRne7dv1lSXe+6Zlr39pMyglP4WU9V4
r+j2eyvT47sGON/WPQNqfhJmTl6VkyFux/S7GhBIwX7ehwYkoqFHdKZSm+2EKW6YQg4futNfFN2i
UdU79GXhGzte/ieYW70wpbZHKH4W+hb60r0Ao2tzCQ0zKDYYMRcTVEdRuf4I2DhYDfhcLAzkVkmR
LsD7TnHPdPX2X84jHnDdg1ivm8+dGUUqM0AcBIMffnniX7FcWloiFieKvLnBDw4d/4vqM3cxNcez
TutPMJ1N1/xWK0vopTQYKyGo2spZHqzZH8HZ8JMuQUWfwiw7iiprhKSm5LPfbdMQw+XxkQkJpZcG
YbKeYIAW9mxantmMXt3TZ66feztBESyLuFBWcTovI3Jfiu0Qf1M9iyWO4yZ/thFAE5miTMNJwTly
D7bv/7s9itbuOmCP2LZ1LBruG2MonyooorBiCaum4cjNu1jIp1PFjw/ImAyixW7+I8Zg5f7I32bB
1WdgjTcdyW1OA+AsXYckuRuT/e9EodUf7Ikziz1ytbBscJIpYlPisZkG8UpvTucR60CbxtWGZJjb
DwOwpx7lFBwf74ERvHYvRKwbMpg9i42VVMeT7/jNUhyfnfSk0wIJRtAQ9xD+SMx8tluTvBKTv4Rm
219znndOAzqyjZMq3L4YI24yTlvnZDWoECKqNwq2TBjCIZc7IN1zU77KvDf5FR3edx4JLokRf6JY
25n5fpFCGamlmwp9Nxe3iYah2TsG0doPxu8XUqofpl/D8oH6Fepaho4NXXm6VExoxvh7TX5h6JzN
ucenm3RpoERsUMpI7P5Ff/GNI4U4Yk9eTmITcBtJ+g8SRVM52VI3Ei6v6rEsccwS4HuFnDon2IfR
c5ftWCUfw5qbVQQFP2x3wAuPvU9UxzrucCrZu3zWBJZqjyFhfb/TJOp1/yX51aX1wVp+XiATDOxI
VRY1I2RM2MJfB0nOofKtY2tCYdseM4cprCclxTTXHnBG9vkPJuhFZc5wbsrXXCkEWyI42tdhTAOG
JuJTyXmsn7klsm8fkc11fmOGV40SueY+xvO12Bq0g8Vic8r7VLOiBtmxVwCh88IFT3zh2Xxtg6Bd
LGyZimHkbjz3PJRRGqMvZ6964Qf5RPd4p8uLmhvEnse3MghxfOerL+ZAMfcixWzPEyuxrIVMRZ7E
8Gci4w4lDE5H68h8qHCNjlQ6Qwvb/JtzepMNHALowbeCBZoynJ92fboZb7OsUYkbA5fFFw+pdW+o
Pyq0RRWPdpCDgS+q64t6fCp72FpZ5heIKqJdN6ocmhiZqsaB/vdpQG4eJpfCw7G83Ib+UMZpzJgJ
sv7gAssMjCMkV23Qhw88BqKqw593s64jF+HslLP3pwdhsXVb74kFSIO3PkBWl4i4dkkA3V2NDA08
qHYZbiClLEDZkvs9IY9Hb0U+yjwOo+uDWV3xHUkNRK2Ov/8nbedt1qiduAu4w5sHJBH3cF5fvw8l
kogTXIj3ahCLNam7EpLfCqMhJ2shpqrDQhS0RCloKdLHeOHKrZI5GF86rJDMQkIL1I3alWIUrKAO
BlX27PG7H80AAKcGJbEMtxVwa2Paq3XPbPljYxO5zag9Kt7mHqVIkK7ZCUrwXw+KtcFml7cG02Ue
2QY1VrOr2PiRa1rttdObjZ88lVrlUP3orFZf/NqYOtszmvAg+h9pAiIF73GqaLjmIWyNMgmGrGYI
Z6JtxqinPCkuR9/0RWcxdiPL+rHdiXgXVVDwIY394wBPDElbtxfAerUAQ/Q6EcYhJiWT6NVWTXgr
mnB50Ui5EwSMrULRXlOGtGFE6k0APPhRgPFTWh2YcePufr4HagaJks8pRW8MTsmq3ytmrsIaKVfH
qh1Mi6jWis39JO3p6sdrYFiQvORc2P501RZS17nat7Iz4hISNm/cruK0KGnlU1w/doIt+8X/Mfua
kSqkHEbC+bKaDkZGkCOcxh+etq8Txw6eAYPSObGw3b8h8i8fCUjFOn1g0H/NKPSB2s4p5TpCk9JH
+3tLMhqRRjER4sEsLzCNLiidyBaZvweVEr3Xi5Ytc0D54vUQObtuLwRKu+HqjVUV9jvRyYAtFO2L
gMQe9uE9lIa2RLZJ3aeRAlLvwNDiMnVrtkWVO97/SWedD8Jx4VROdXV24ODLRzBkZ+i1+2u1ifZW
uQkjVBaevHyQqWJqIjJFKHdw1jyEx3JMQW72f5VSuzqMaWvX4D8f++bh5hbu7nFBoGULZ6WMQege
Dmv/HfwDOrLRdX8TnsSRWguexK1NonKKu4ux/J2OZhGMsYRaHta405Th4lCSPFUQ975lRJGbyDTs
rjlevXi/TsTajMq6OiTUVfNzGRXP6rhKKsUx0gmzcQaLCXcYfj11h4sP7V39DKytHLaiCQw4toNk
4vJMgxFT7BvtoqLgZAHnY1/FLxdiybnIawHcBBvyII/MSd08uR86uP6bvchRi+lbttZ2MddJ6Ens
BawkstAYOcmLl2mBYpwY97qpQygud7Q6pxCVtD9kTqMaE+yDQHNPHcpANu1T0init3BKdI6CvV1h
qrdXCUhGelUp/QQIGISePB+Sie7xxck49OLzuyQZ1yiPG8OIHhg0hlTebbbabUiUaNPpzwhNUbNZ
i092Y2A88Cy+Py7gYaXemtErM6QL44i3zVymmDhCIwh8EfA7ia1ABidpeJ8lCPvYtv71V0A5PBtg
dHTvpWlUkVIMRYx2jxX6tBxx7PwWgiXgBE+LGrQE/oKOm8tI3v91dqp0ecITqqbMVbeX1KcgpkWk
xXAZG/licAe9YBeLSQJ4o1uTvd5z4b50qlWmgCUBlzxm4sPQkmM7y6eq7xhEsHtYfKiMQTewywRG
b2IDrmHXQiCnxYze0kMPQPPfCVo3RyBjhxuky+epsI5Pt9abVg7u8Ffk7+CBQdZrR7IxA7zu4Gkj
4APvqo0nFGdqJUrhLJqYnTL1cjhiGXyPvKXLmXasDE+2yjs5USq0kfz72aErZchSxyQ9iKdZtnz+
KoZFmwA/Wc5IFfQKMBchbwSVGoIJl9+tvbvmBNoOEwp7osyX3wM7Qlnyc85xjXZIYowZIdvrnkd5
DIxOpR6Y8KL26D7vms/R9RYyFTNJ8V3Y1h7oPac4ErVtTQsWjJYcwxS5gTyDCqPZEevzkNJ3HK1f
9M/xnjOwLqw9BWuQ532Ny0wV4Bxh9wiutG9bDk/8cykwkEtJhbzMU5HORxVKdbiYWSXj/xag4du5
L8iA18O+9Gv+OkX+CV3jf9LBA2WeFyuYbEl6NpG/5CPJzX3CWXADOMv/Xb+s/eHjnQQkz1hwxEwh
AqR2h259ITreO4zUcQSTlpvUnQLwGqje/LrMI3cKH0sivk65D3W7eWAxhKFe7cJZjW4WYeQxKxYe
ixakSPCx7p7CHIX2tK0r7dXTMP089CWJOtTcOfrnI3MTxpYj6G1G0z/bi/2QTBFPL5YByQ8wummx
equS4Q+lRL6zl947O4aXBCwQAnMLbCGX1JL8WCBOD36mPAgw4jcDzp9nyUsNI3wcvCTuqlevG4Zy
GR8cO6Pz84hXOQiO4WVBPxRrFabXaFe485FBwT9KQ7PzkDSyll9EfyfE7B+bqbtxeGclfp85tsZm
EfXFsWB3PQt6yeT02scGfpVkeE85NNkFaPfHCS44JjFcn3RShI4g4S4glBpxYRJlSy6/0utXrD1R
p6AL5osH5yKhBZZikXmZtWgkLBeF9dGCevNjQaS99HeB5GMH0jXso4/4YoyCWSZTx3wJhYAeE8FV
UIo/vkd1U2neY2KwO2iY8nZ+DeBMYLg18h0urkZeahUon56aYLPnOwPiRiNmaJ2A02kszKmvOYgA
TobJPBEXwL1PO72gykjji2uO/TypUPfgFwbRATKXkiD7UspmGq246OSpLmoAEF92YXIAnRs1NEFN
b5eIHB1dtqfk6I/JSUAQoy8+JE6b3gjWmyGUq341LWh4klFd/WvnoywxinzcQ9FZJEsTHf4oJlbS
8WSyHUBnyEqGLAd8x8pf49oQINGSOMJTBm1MScC+mSrg3yozpXFgr+Wj8QkWbRgCXeBWhhmLvkY/
ShAWrTr5kjSXjxf+Mkp73LaW/jmptitjO4/9vPXOpUwx5gDvEl7ZFSz6UNnvJdgRTP2clrC9D4DG
IVxPYwDtOqXmqzqrb2BUOb6p6TJB/hxn5NU8tdcHk5F2TrOYAeOLyMvwbzVLWQmohy1K1xglomFu
ZtFc+8TL5Muqgi/K7zswqTGiMR1t6jixbU7odDnHrnn+xIe3k2kAQPa3uC/D8jArdnyw2PpAkfuc
49KjdH4V1rjZ7r50FYE8vxrPbbLwwhtC+mEK6cvuqqQSEbPhw5CIUaVZxXk3kPzYYxOVXrS/n7aU
X+bj3aPNSE/Sxy7p7vkpRX/WyiGKo9QN2rTIChcOFViNl30lJyWzg/5K2pj1RodQXVH34bvk6S1w
OWeZStc5uap5sH/PoorWAv99n0cTSvAPH/QWkMHFw7F9LxX+pZuBlxS/MwyAYHn71eWTvNgO8Pgu
u2iNdwbYBlPJVP/z5TPZCCwWTVx+QqUI4uFeTTAhs2CRNBI1lUkT9MSnjDiLep32QY6iHcZ7LgWc
oQJDFWuVjiyeZk5vjJ3lNJp2QErrZzZ0oL78vwFexjx6QQ6tQr3170Pzs4r/o61UOLPKbHBYgfQo
pAggGnbghNXYzLrDvDaasGrH+g0XsSvyCUm1n/CHi9403umuhv5Fq66BNVZPflaKBUjz2ChK8Vat
JUSprgOHRdkCHTWCa2beKGrGfxrQ6MNKe9YthXsqVTQyDR4YjgQV3wKR07YKcGxZ+K+zjrP8Ef7r
iIAkPKXoXDIt1mZeiHQlrqO5+3GiC7C/BzkTdypyTQv/b9eHMeTY/D4hcimIrnaO4x0UHnYCojjM
6JRFNJ8Xhanksa1t6Eh81+b4uGYxd1xAfbJOjBB23Fwn/XH6p4HT5DSCxHEAGjycHbk2FUAHMBU2
vUObRyHzZN+3viI8wWSYqlsA2JlWCDzKhc88eLv5N/kYrxNTPd1/pdMwZvilNMXnwhqvFQCsMFUg
Riw7txPwJdoe4I6u+iRQi7aOV6jbU8jbPHj/KdQeiMC9DoQwF5JJFkJv0/BKT7oPvqITeBg9w0fJ
AneYRC2hrWmrhVbT9/rtYRp7FGtuyYQXk3FIQLVARSh2ta53bY0vciEnmme7m43UgZN8s06xuJJj
RHY4MxVc4s5N3ATZgMa7WsxUCVNe6LAlCPPmBVBnexWKMXOECJaDyDoQMpccz8TKZXXK/xWkzgsh
RaR9BgBgF/2xzhhpiwAb4oC2FTr7P7e/JnNVD0aCD/ZEkSEemTpNxDfPK5hk/4p9aeO8D6Dh9fo5
wzaIo+/ZlKNTj6hDZZl855O/Gol8/ziGniRAVe8XJDJ6oj+xFfSAZR+EWhEGfok81uRCCQSoSo+i
Yg64z2pbK/uWrDYH9F6KFx62FtqdVZLc75mU/igtxXMsD5/0Lous02Lhf0WFYQHhKBuXxTkdYHHZ
pfFGXzUXZQUZtyyaa6DQicd7kNA1QX00n+UPJrgbgsNVXgmKrjEraR2DSQpxe68fn7R/8GyzPcVK
7A7QZGSUvWtgU9OeltCFfFTAtNnJ5uj6WylW12V6ANXsDaFNJXILB4wdvN9YliJ1DWMz6Fec/5vk
riNZ3sEPTlf8KhP/ZPRQ0QebIJWtr0zzHC5jmtCVdD0jDeR3wdj0IFCHOIbKEBoNRXla0SdE6EPw
uQ9ShuK3catNgM1LL09Saxl5sQtfIcAKVnmnXy8LY5RqHsQiWyrpYhpwTbMIUVVg3nXisUeXYEWu
2jZNU2/XcjKTCyAUoqckkULF8nCow1ACBbDJQcaM216kc1xDw4Tb94+hxFdtvqYmwLx2k+WbZJB5
S306iF6hv0+Fbxks4QQMv/Yi/0fEb/f6CTjNff5pgAMImCZNyubKUe52d7t8QGb6NiToxUxbZUW6
R/16AGe0r4HrlTDZ+ebIkdMMdegN3SrRpHxCAkgR9dVosEUmOqyGfjdVnOjI46UClU+2lZp5bFRv
GLPiGmc5nlF7US1x+v6tGkfRZHD69ikjEDfsjHfJNBIkeglN8aMjXoXSeWj3OTG59AMTMQBksZzo
ewcrBqt+EvEqf5SxvDwTTAxjNTbumbWb+vAhqhbTCnH/1qDeCocmSZ9+U0yKYu+f53AhZ4d2Onsg
NWNJO+uErWsMq0YJa5Or9IwLobeEPXrx4H78IT+LeKsv0krzf4o7p0DTtIh5jWfZb4zd4ehRXBwK
6Zu5EQJw+AkFxW0FfqgeleTB7k0g5UoVz7jvefMsqWvah0Jt0FIE7zUXi2mn+/8bW2IDuUJpkklr
nr1ssn3GCX5ulayNPFbQZVhQCK0wvQ7zXoPiqtA2BSmn4g2Na9+CCqq7f2mixQAAwu19hW0Fegpi
Y5+/5/GT2ie8H37BxgEPcZMAVcVCzaOqS7aOEoVUpjfVxLZabm3fmuy4qWbpmCzxGIKogWXnI9d0
Ry/YAh7WkfG8VgBUTm+qAw8aFOl/pP/9MWkxbZZsdpV8PUgcSwBs07TeDLT+aE24v+ue8NNK6SlP
XS2cOQvkXAiLFok5746GuCPIy6Ai4nQsBqcFYzsR51g+8jixWkOMgJGwHHhYmETJn9Jz6sSQKCmW
DRE2hxeu2d4QOX3WUXXEmEXfzCsvzziB2Xq2c8mcfa9088OB9oTgRwSAlJQQ5eFtQs8iS7hPE4aC
cFxscoLuiB8uTPDY+a1Qnr+nRzMlhCz/jJULA2QCgT/pM8dkeF2lYcQR/pyR5YmZgLLd/tmSlWSW
BLwtY23+u6e8Vc4clV0JwPsH4MZda+zkwQjZlegSzzogtIZtceSZHswvyWqeUmRl+3OWrFCAsMm7
to31xJ+0pFrDqCRpfG3SENxQG2nNs0BNGhCF1T4FOGQuv+l2YRzMbJTvKEeXNZMVXcYBrEN0m7Wy
vLjNccP3sK3x68IAY9QV61REFRCSmOJzT54riFHXqYnMUvzJZq781DEEtBLMunBG3vpgZd1vFkek
otoxLwrNe70GjQcSUvK0TXN/b8FCOln0rJfMzvU7pBT5ZVv73xD4eaZeys8FlXxDlEL1iNeeOwk6
AVmDFKxU4ItmHBU6mkHW9UzDoe1FvrlFttNVuKeSWVrt16OVC+7JuS38q6vv3jXutsC74izO6zA7
m4d/ytkoGeLr8PcEWx6VtCGl+CoANhXWyRMuYodnO9Z2kbt6o2kN4zKCN7W5pN/uhj5oOv4ohEau
KiVtjQXr0mpi3k3qvGgIHhtExMCnVlD0dnSgFvkbtMtvizHiLwmTTl+4bALY8vdUVdMf7T5IA0tu
/MvO8A8NmgKjhjsMMwYKOA2N9zcf+lUl04cYuf2dtcHr3YJFKOFbftpiBrFHc2xgZ2u9lHe5qkhi
hhbSWJNniafWka0FZpo73jc+GMJa8DU/IkfH6ma5Wgea1eFtH0oJht80FjSHZjfluQbvItf/3l+f
CUTPCN+MKNCGgfqvi4Dr7aY4vv2fOj7payix0RWuS6oanHUHngYnDVtS5lEA42jXl+gwFpPzyCOs
+1VymTXNDzZJ+VLYw1HqfiUgFmPqj9a+FdI1e3a0oGrqPUznt68lRFNgsSss3mkbgP3l4r739FVR
Q80eE9ZBPKWd2ZcoC5EpE2Tfo/lmi8+R/NAx/ASpxbWAg14UHUJqgwHJIQisIuVxtKg5GasgIoZB
tcC5y3i79HC1OJEi8x4BCUXSrbkvOIXFxr5QTNdcPpWMpUl6bvxIbvZFEMgSiY6s1zFLdASOhxrz
J7PIhuN6f2mY4RVRmZTP03qBP222Zz2cVOycS8XcvKd7/D0eIxbxAwysb6CN0BroKcISJ67AWw+g
vLFFPZ0T1/DzojhOs5EMBENpuztZS+1ZkOpPUPVVG8fjp6Q+ek6WqCPy02ifRPTJ6gfBBns0faET
L9SAxkn8rm7N28CmjrHQev4qT7bY5u4cdADR42lwJIfdGozAIStGjG+5UMleRPyEq+UQA8V+8B6h
ljOMj1Va/J+yOdN1szJaLBhSv2UAl2SZitVjA9NybfJFB90SoZL3rbndSshInuAhJkUzVcAoKeVc
lVLQ8AWbx/ye0CxGAwbn6v14POQPzI8dEclzR6A79HXhYFMJQA8F0HH1gWfgGD29R0r4aPDi0p+u
YmuuscoRGv9PktWo3HtnCDn+0dFzPLoYVuwhQ8ruCjsjL5NWG8+ze8YyhNkclQOLNXbg5IpiipME
5XYiA7LuX3CT6QwvPA1y/73bj11b0ExVyvh9tUIaA5kBSLaUc+Cq3gmyz8wp/x6x2bAoS0z8XAvp
gtdAcqaI0UsJcQq1vml/R84OXn0gMM6TBfUkuaaabHXzjYX7WwSe3gXZrAGV7VNJsRt1jcxn9LWM
SrKodVQum/gqRW6JRHCKiWAfVbcEYJoETItddnsDfysnsJ1GcJfO9Wb6SOLPceKK3x1/XXwWmz0v
uUE4b584GCJiLuz9QruQXJkSLQ5Ch0DFeskgp3jxFwp5dEV2zw+bKonh6BB2vECk3iNa4j3fdWie
oYYIoXuIznC8Lnc4keuxA4O/JolMjJgMmweNZctcHIVJEanRYaXeJJbuPOaL6uIyWGQFyuzoZ0hk
izjV9qLsGQpmg7WWQ+5mogdyHlJY7FO4kJDlTz2FOA7oOsdB+c9QRS24gDaY8oVnp3Eh5HE6N66B
gQHsUaGf+mqZUjNrbApXgcQKi0XeWIEfe9iuvb214g06SCmEK18PFxMG1LGNL0X92xt+Dx1oAT4L
RXvJYUGbDq0ZpDaNtoGOOBSvmqlZ9Tap/+8cZuC5FqSGgFjvwj+eSpdumNlj32vCejgcD591a2Lr
oaqP0RknZMv2jrdip5CHE01VP8lOzdOAO2oaUCSq/hT78TZmiykKItVlEOls7Cy6okupldW/EZ18
udOJVHNAWVaXnGr636Sgpo+SNNyVOiNu4OmJ9mpcwZzh7gc4AavGNuppEQ/1swYXYpm0HLZhHVE5
e/U+V2tSfzgWQCI7LP6gd0CTZuOYKdOOJFHy2JwX8H4rix3Tlc9a0axoYPfRfuwbqveDNHVFfY0Y
gtM1fNhSxNwIyLai/Mg+8MGJBziGMJJnCKAA7PiUHvMpZboWo7i+7PYmtngPlDy7ugSvnN41bdwl
2VGOdLp+WamlWWU7VhWzQYr9cMPgy/4NWyXedbu2d/fBTPw2mPCoac2uh2SF9xF+p/45MN+2tCl+
6wiWG2nn+DEsYlNEz9TkxlN+UyZuBZPIztfetwl2gBECL1pNS6v06STcs49CXutngL1fcPC1869d
OFboi2ioGecZ6QSGLZy9DRD879VHVue5l1fz8JaXM0c/JH84XRqwnES3jXUa5FWHozY5D8U3DPTs
rltm6OyGJfAmaRSnnFG7GLzwCJJ483xRRVAgUnQ1mR3yGp2GoRtH2zHgZMdC3nKwX1XJkHcYE9Ma
3AyGM2qWJap6zbGMEvlE7ZkdLDtQsRezzFMLb8y6UEHU0TNu/9Pl14WuERHfc2cpVJTQ478fCRcr
FHv/ixbQvmcP9RnpZpm1mUKayY0Tms03i1BHSHJwU8FOMgbxzVb/e1OeNSR63fPbf57dVQc6Dnlf
Rb9kHDfatOSqi1Yxg6Msnu8g/E68ovYQl61KNj6CTMenK8jh3HC0A2mMiNXlGNaa4p61Qqj4qlub
VfNO78emMgQIvynuyZFuTgsd9QC+9zYQaH1usyFD2lKX7EB7PNrJkEhGKxedjmM6mRa3wunxnE/A
j6o0mxuJ16abMX41544M5Jc/buKpzWv2KcZ/6LTAMnuLBK0IDpusSMwq/CflhZF9/pdu14pzO8SA
gSLj5Ns39sXXRmZwU8H6BV6Mp3kKn1mi9D84wJN/4ouGgBS2CGlceonUaW4MB3Mw28xj3RKG9jm1
KumSKCmG/T5H1MEhvby0fmUF4izGHBLgX/oyPbH3YRC4z4YwVR/dqKgOG9GIp4cqQ8E02eBPiaad
HEF72lVoLc7p37PAOvQyNK4iM6mP9lHUzqhsWw9MtSJsCgK/47W8TxJz0cgP9lhyzuV//rnU12Iz
uOzO7Wp7HLmsFVVKQ140mQ9+J7CuqNRTpjYFbpa+UBbwAXFTmPt5Hcf11zQCnTypjX2+BtA+ci4e
RKmljMs1PLPdF1m3Toh9vyeme3dCdTgvXkc7DTgH8DXy3TErJSBLL2ww+IOCtKVmXsKWR+cMHK6r
kDePiv61yXHjgbOJ7LxzvNUwWAXfOiAmgUJqsKjriVW+B55pdhfHvbjh+FbhpNTEHQcN5TCASn3W
zNiO/Y0qHQ8FEP1bZ3A1/qI+F58X2xjPDn371yf5ZItSaonnuD4883nbd/hqUOkDvVfrlS1Dk/h2
TYY4USC87rExI6Wn+nt1EZUPE219XXs+a1tmCZaAXt3lIFfDzPnromENQr3UiDm7d8Ypu+9chCFY
CT72qD9E5HR0N0woUpocyE3GEMbRxQ9BSn+eeRlIphN5VHQ0RinpDzIKCcPvbQNjgtznIIZu4wzF
EJ277HU8606GFql6OanZA9ZgmajI0UpuDww9ioRckP/lyadpCpNOP7bY9ExvKHOAF4vtST+e1oCc
xsJOeHFI3Vk+MPKUof2aOcjsbromokPdjwAkAmMvTGNyH30Bf6Mkvh8P+ZNpVvHKDXFG+D/CQOyJ
Jyg12/3bdX8VTUNSgQdW4TMtqleB6++IBalBA67qATY/s0seoZku1oXSlVaE4Jwt1elXmlQHUN2c
QwdJO0RolaXuuDQDzKpv8UNdKSpIKWJcXBP9zHnCA/aoQhQuNG3bX3nVo8uXhd6ytNEE5BxfO+45
G9ROSgZB3GoSKhuMLJrnp4REuzcKmaMx4+lYAtRmpC99Z8fXfWhibUJfkyMoDp7gEvktgMspCe5s
/y5MvolGfs8CFeKv8bb3TzwE6WCB4wHdE7A1x+gA7eQYyEHd9SZ69Sfo+WwIQSnwA2b5R/GiJfv0
HsBQaz/9uoZZDerNE0DX+U2KkYFMg6KiAeofS8//H4eeAwXznMZETbJzK/C10aMWEWdP8ywzeEob
NpCLVr/7E5Hp7Hepw5DME+qaVfYsWEXUnXpx9z3zDwrAOwccFqpq/+vVVhdHxIiB5hfeu+E0vvMS
Ry8ABXxh01xSQOysGWR/Yo0TzwyzLYbIZsytn2Tsg9u4WKW9aM6Ffkjev2qsDhp7Qw1H3xCHaD4L
FHlIJuZugTjRbQf3izyMZZK9/wdQ7ZeObrN4lMMZXTs/oz3/4jB64PeQOKVFNDZs94hdVxw+FQ+t
i3u6inoeyvqxUiCnDIKNcHIhqiAR1AWQG1kO5xcGpytp1rvNYKSF1JG+3EiWrMtL2ozfKGMO4GbR
X9QkXu9PMs9+aKiBXYnsKJSArz880xb2nKHtPf2C4sI6Om/QmmtJbliPSZmdIKLVncuCICRAm22U
wKVtUf+ErmLXba/M47X+oj4xNTIlScWWp5IraSJDPxjPZ5ZiayO6C/UQiJt5TMQwuI5JQ7eo2Mn9
EjAGOvMw0Bbh0MFQhTBj8UvJFqwnvGrXWyt9DOKORIrZdAGZH7CTMs+yvzxgeF1jblDytqvWwEtJ
3tE0NwuuuCKqeUNcztpMgRQwmy0RCSKtV5zcir9a/XQTuWTljiILFuz7N/i/nSwGJcYx+nUH/dbf
GnWS3nfkUG5sMiZLkZEeQdfDehIoakOnXuf3qOrXCb/wQqrt67g0mxA1SsRn1AyYqERFzc8FTbwa
L/0oIbMKop+Lb0MIy2d9VoW9MdmDMdA8kHjdmrywQDST+0T3z53gVzT0rDX43dyjMsYJPBgxD9ye
9GIOXfXSu481zDBKvBhEb9lMXc42OLc/XuA/divm3U0EYbb6odJqplBSa3xjtbPlTORV3YAqk+K5
zUiAO05U50mAatm+xBQQNOyEQKJscXj1VhDU0H41+cW/qF94iTcfT5UQmaAjd1HPS2JnKWT0W4eG
yVaStJHw571+5FCrsaySj1PEuLjsqfQCt8dPrhTEA4HDBe4HsS3kKxkcWCtfCLg+Rgf2TKQpWT/d
te0FDqYj/IQHD22B2Lg6szvYnwdUODzlVz/jIZAeGWdg8W6j6EMLsOW98KxZota1oSGdPwMnQ+lg
ceC/FNeqodGJuvUemOdHnhBmlNlIGaFYXIv/cM1KoQuTqN42BK/MBSGpp8mzrpn93UmySQQepqaK
xC4sk+kosJMcn4NfgUq6nVYb3hXg/nM1UeTBf2jZr3Ncqyt3A1hhLjfV5iPJvWBLZ3WBMXtVPT7t
8hnhxg32MBLs9zyh7TvUs+B4rNjTnqdiyUHf5FqD6klXAWpXXbPzUzH895Ixb++GRsnjYh9hhopD
iL6DsQnsuUNzsNsJPauit/mmSIvkdYONsJuiwzPNh5l2aua+YqYjT0CM1ZnGqg9f+5FEP4tQY1Uu
Tcf+os93EVY/Y56Qv5YXigGLw3CSuNuVMhJWzqIqvDqLyk+/Vv09bcxjzgUg0L/1Ke1LWrCM0rYU
91TGXruuR7on0KjXtq28Sc5deybHQBIjHLz9mzLL5TbjOmHoBF/JYwshlKxTJRHtfX0uLbHmHPXg
11BEtPtD8M/lzQSdMQpsx5r92s0htFFGbAHeUTtA5lcHJFlfySSsOnMCPK8fDI81U3jBJZssxsEJ
t5PaR8u0kpp83WSALfQiZATJT9Sd/rLQPz+O4/LqRePJIA7aY2sIo2jkp5O06uz6EroCqiZoD/xA
i1wPcM6cVs++Q9J7UAeFQnHm5fsYUJE4aQmyMDh5/FYSiGcXPKg8L26yXKGXYQGK/3OQuP3xHCXI
HzZEfLRXr79bHjncihkwki6j8AfEjqM3oDYrVGY5KBK05QMBPybbMiQ+pye/1vGcfRXUsWJkHxtr
zRpB0+eQmy6v3MD0MGyAlQyzaaME9cjD2Wdk3isWB0SB6dA/pL1k4K4vanVXxxqeD36yGadvC2s/
UYxbqUKesdBBEBuGeWblOKeUyVR6Qy2wZRkmOBmY541vB3OJ9XPDwLeZA4wzj959+2CM1MeD6PEo
2fF3PqfpHWCUr3YLmnPmxIdc0RIjMpRuFUcgjYgHT/6RkRvV1UBjevrSFgR53xUFlU3XJ7oGSllu
77vgwRvS3ITcDZzKFCOP4SlArL26vNALkHL2Bpg5h/EStepB2eIKTDo4bbqbl/HSCCUiUr6c1NIl
FwmoxcN6rBoPYj9uZZmTe388yZtfwQ3vu1EStc5AaOfJYIImfVDUo/cD5CCIGudJLt9+cWCx7mlZ
H8neWq7n4HLxn4+Zy194clhahRlq9acKl+eFXqwp/UcIWWLO/1HuPHv2/8muuAbUnovb3Cq8Im5I
F8l0UmDw+H46VjVL+VEB7i+4aXZS24Xot5tNYfPvuaUY1HlTU3cf0jwG/JH3WRvt/ZczzCaCFQUW
C/FfNQw12suedFgsrYVtPy1PFKgDrj6g6lBYiC/XhUOP6mld5uRrJNo6g2Bf00k0XzsOWKurWSH9
cUqmKalavwnXIbn/AKmJnWr/bWAxJ9kOSMRa/WRKOWO75hVPpV1ujkRrWPGmSW2+gvGQrHHmGoYT
Kn5URpvQUAgYAs1IIxN78sSOYAN54IoNAC1LJ1CA4Hktjk5f5ajVNqnRzQLRfrxzv52NmQ3omf32
30hID6RDtqszEAUI7FCGaYEBC2X7J/da6ChQiGxGcGXclpVJkKE4hisvM0qWC+iHVaXM1uC6QEvM
rRMREUbtmjN2gPn9H5pvvaEjVSR5V8uW8GoKx6jM94rcYz2tNy6QmSugWDswaz1uIiWnttWOsX5M
lsmn9RYnCF0SFv9fbcerlVuJG8PwpoAhpWOZY/jqVRc0hehlKziKNg9U6mdRxohIxRybUbaXGIPt
B5TtWZvVdO0pZ0e9+TvE1vQOC/lYquruaxFNq2AZ+7gsETO3PaCNROl9ZJbSck+YsxeQKvHlkwMh
Cv8SlF4MFF4bVGjyiLg0wZtQPrR1MWfJrfxukIdGiV2GhbaFVpxexFqems3GvgfuFoRGa9WOhIY7
1jIiLAhwCpWdr53I733wf2Z4XlK52E3khhEG5SCtfeHoAHdQvWkJ9/e2JRgAgD0ofvhDmQI+mSB8
2D86nRZNu2L0FVI1DvlJT46dvEj9ctxYVVgjPjQ8r1bCBu6VBFszY1FuE6UE5xM686jwKjPHe43E
D6538jxzQh2oTIQ3apYbn8YSIfTCw8+C7PZhLbVsRNAjMKTWIJakXdU3bOMp6ZxxYTV8MThqH7IT
iSGdxGFiV7nPN1xXpKLl+CBYc+gl0wav7nMzYyH58D7a0bRmFg2X7AJZAiIMvmFJC0wo1O8ww4MB
vWvqL+FmI569OdMWdYp5hkPFkBfoTzAnDnYow7xsLhFG+tfXM8DmbheBM0c5o8YkZUw5a0g3BVeW
1+M03or3sqAq77gDe+P9RCUW8gV5p3I+rbuLPooi+TAMWq/2sEVOIus2C3vELEEGQ+fpdswTK1Ok
366w+fs2pBu5DE9UaCDl42Ry8TU5u5rE4cE4BtQs5+vdsMOXvc2jLJxK7BGWq8f4D3gNKdZC8cpl
Jo4vGTYJeiBygPf7SfrJAd+O0DBulcSpsCqcXrq3OF2vTbm/EEGoMuxxTMca+YprCpXwWjk7IdVS
CqQNbLz2BTu2jCFZzIfm62T9yuH/C3YTydd4JHbHRoaBxm45M4j7IzX/qS4NsYcPi3+axEc0X81T
29PUTYru7sNi6QV2uyxhJaURrA291qvZ0qmq4m0Xq/QAUGd62zrUTzAWVXgL86eu7mttC9+N2GzY
wRn3Wnsr5ojAGwG3HfGhE8DVsQhjMLMqUCYlsAaBQDAjGEKxhVlm3jQDm7WCwYqGOO6I6zCWP4zI
0YP8eVOhXMArOfaVNnMUvwVlSSgSj2rn7zzM0EBkiwfepVgYGrzDoLsNIsFoYeVGYWHdf25qDAiL
/QH6iQ/WjUqLA6AbeNfQQP1zectIYV8e2FwOHOZTCMpot4iJTtMwhumEJZejh76levLLnfGlTKjY
PnxnBIGNfDOyGVetMt3mInqGGUzugSkQnWCm6lNZU1uSmnljAGX4SiGA6XS/4xwHKELTEZ7pYlAe
7EELGFkuWJgldesK8j6JZMKLNatrB1INqfGdkEWmx/MH7kJzP3nLewkZxFxGDrGWSNR6pVnqV0DF
4UjlCIREvSpnn49IR4ywz/taHXBtdMsN3V0TAzjJ61tcZuAGJhDHyVfXfyN0hiWRhUr2vAOjXs6A
QAsA2o02xZCBwq/XsL+/um/LUb6n7J8r4Rdqzj1JbIEO2etb/6UHLgsM9q58/lDuN6vQNpi2So9i
Q3zvyUIlQijQroJBBczoDtJjPustJUvOahZOCvlzk5mOGEYKLKFQGZeVClSEEEqBhLJb43nwdnqw
AuJHh0mNOstn5VWrx70p2zLKvY2j0oIcxB7NF9JpF/k3QifIiiNRdG0i5iHf9GR2YzGwPpmndBpO
f/jKfR2rf9KOhwIjaPS91R/7s+3YfGLqBkikRZy7LSe4DLNqXdNX9TjrH6Tw3p+8TInHYNrOJAw0
ymHmNgvVtPg1hygAlXob9cAl5vrvP4GdUJDz0t4JAAtlXgaCEgtkb68Ml+lfB+RNPPuKem369Jd+
DbTu9Lmecw9m70VZQbKYT2IgHNsw4BYY/nJ6FzXc7ZCzrKLJ0hhWn6BymP6BpPqI+UEe2l7ZEua4
RKYcarD1Xkrp5/9FPWJtXPhxRAy9H9TrySSNDaAlN1gxckdZj6yoo8d6lc0jTwdccv4OUzVDuNrz
JqV+wyMZXNp6Ux0iQn9Stqfd8pmN51JjYsjfjRGqxhOV+xJWA2zyVr+nKgv9a4aJxBJsLjEYE9DD
ia2iBRsszCbrPSkE0MzioBGbFOzgQCSj5le69MkvwfX26FIqD2/Q+D69h0UjUNS+5x9W8ylrHkpl
Ja2TFaSSs2KRyYUmkQ5Vf1NsF3+WlpPyPNctidYbKN7X9HaT1G5HhHZt36LHxj0Fm6DRFDRhbmAk
NRHFKx6rFZoUowtT8YKEtqxYAmns/A2A/g8rfQ31KFqETwZz90dfYUDQa+dA966nbmDkD1Zm/lkp
V++s+FyCM25t22RMcxUGX3J/P/xM4/Bpfzb+XLALnfWm5rKTWkhxH21a6UHxLfZsRkTtmu7+SfXE
qxSOaIgof1LuxRMe+UANBfF298BKXAiwLobw7guGoZz5HCI3L7YpMRi39rRZVuc1UO1orD3/wtta
gcgsrTmorKjISdhOnUm6Xzc2gdCYF2vJ7OQujjUtZx2UpQ/OyFSA9MttThhloodsVTFSYbpNrdQ2
fy1Nq1k0vKYFUKxe43KVgb12za3XrGoGO4n2YCtZidb58VgV9JOPorSIG392VhLHJEmURmhm1Cmv
7rTcOEzynLH9zq9YaBi+kkyRY74u+8whRKBfVpEZRCyUxl7a3Z48QmVEVlE/izs8OcbgX6yu413L
O3+Xyrkn03jLaDjgNhOsB5bAs529iiiZmWt4NuW3cr3cHVpyI0tU55HOaHeH6WY4ayYTVB7guBo+
T00N+dtTHKfsHOzSIpduapDR2YjWYot8EsavhM6XBYBu0jNaag9U2Mi5uIrPUJ41OKutrMXANRnD
Sif9T++F1+26xRqmAQ+ZBPqVyJ4wHY0gu3HKKWA1wBr3niy+HAvLMapYvvrXbPBQZqthi9aRy690
8FwfI57h8XLpdquzRigxgl9BuXKj3AfNpXdZWbfYX4m1hYBzVCaSsRQW+pYvgTh8bGSY8j6V+8O1
85BilKehrPtgVXutah8Dw7p4whMhIeA+sw7ej6F1O/0p85x8XqpN2VOc842fYQ/ZQw/Sof6rtgcM
Ti41aQ9y7e3NCXGLZrsXi2RU5uvCnITlB9qBVhB6y9qP0lCpJFx9T7UlSyRx3vASpNeunt+9VwYO
oESCF1qDWDnskmpw4phqnVVC+ZcHSSzycFhUs6qOa7MeKlzBrLog1uklmvfKXFiVne8Et5K5+gPx
iqes4nA6kGfqmvpcjmQCK9Qm8wmmWVECCJdMEfq3jTbWwntD3miHBE9Q+wHHqTyFrLRYpla7DTSL
19B99+ZtTOKqfHNxXS9WFD3zRpVgUuNhjcZKbmDh1iOffV1OcCq9vbgIVW7OGWq0ErIheQre25mM
lpE+292T0Atje3jYNb9TBgipjfwBfqdc6JawoIOeLQoIVgHahsTh6FvVt7ZAp0KHJLS+f+PPkA0h
a9aTF0wcMD0Z6U3RwSuB1Ke5jhikBxWAMAwQyQWTZJEVRaht8dM17AAojWqe8KyiiUopbIKeCuIZ
5RonW6j4japnlmSu8wAxzWmivqcVdwerueorOCKjauJ+Ay2QCqAcKVHLD1WbuR7ACohNrCIKz8hb
ewj6nGwWdtTKqEEeD4LL/yUSInFwldOQlIzYevSgYTcqwhrHzu4uq4QKHpjSrnPsCa3B3YIDnlE7
sze+ARIQeS2Q/jp1t8Rj5iUDNds83A/I5Ni8BgDNTXVb2SG3ViLA+jrCf74R9XC8MUQLI3WjN3zH
Tm0dzta8Rt+Uzmh9eNpLIe6mN1qjMa19LuQSe2ywZxoNht692wit/EwOO9EA4U9yzO55MHbHo5Mp
L1tJ0rqSIOL5BwmvYaJvQJjJH4+NnwhDt5xvUkDvC91cI4aCZPcDyrhsDBPkHivq0W3kEAgKFB07
LEPQbOr532dpLbZQh9+sCfHOafdR/nDDeYfxTYk4LfslQ3AoTcYIdTgzhrXent4gZJqrUM/KGjF9
hPGaCe7hR/lfm7im/O33Sa29GrjBBYJua+1+oTgdEUH7fT4bsUTSJCzkLu3p13xVYTi7vny+47RF
yyYvnn0CkRplrUMH3BRngZxdJZ8Y7xNDTGvk5rRaaOAe6yk71M4VUXeJwo63DAx32TYu20bQ+kXO
udczucYvI4AtgjDt8B56crE+OE7VskbyFU2QB/yqn06OQuUKF+1UDJhkGOYAGJR/vur+qRJLHEeL
gMz7YsOR8epyoxf5hm5AdykCUSpFAWhpGVRZPZfgC7ptfcfyUPtLTUgaineECYvFjmsN37TEB5Dx
UKj/YOOtEcYFBM3Mytg8BGRxNbC9nlMj+eIJTywHnzBimCcHD/xjPwquuNENSYYfrTGBPNLLOaQ8
M1B6wntQE5TTgfj0iUzW56R6zwlv7t3Lalta9H2znj9Rc66Sn7Bthjf03V4DwVQk5Q+BAz/Kb5en
H/DzInxeDIl7y2XV0NQutbDodTM67gUA1dQtnC39NlELkr37n8Mnq1aEDsWRlp/VRtCyYLIAAVPr
bP3Tq8GMgRf/FasOV4HLedRoG2ZBqPIPVICE3RInVNQDRrBVKTwn7WkLqgG32b64WzERAvjZicYs
j58yOUjKd0qDPPoiLtys9upYdMrKNYMYrpLgKjo7uiwBQ8U7hfGFny9xkai6YkXCnA+5hHgXU/U1
49bVOfWoMgmtVSHZiVS64X1fhKUUikjnDzScb8GNyz1G/lXTQTL2PtUv12kkd5E3PdeNCxl24Itl
cOZybsCBmDzBmebQjV8bxvmKfGMdKBuFTpV/9jNQMeaH/S7RKuIOC+RaCYfiRgI6SdjNIZ/y2g4d
jVK7R7DZ2jvz/79oK0BF/yCtIsPm40EAhO+4au7c7fLRbLhFD1tlrOQ174X/YGGAvxTS0Nd2Hj4L
21fAPaQi7gbark4BZE5AIru0dqtOEWtjzujeXGEDXc5lYzrxl1AqIqcOikb3jabrEO93SEN+aWy1
HmcsSHMsDIuuIhk1tby13pnO0uzZUFS2/8n80YdNiaRRYjYQrh3Go7IdWPV+gp6r7rGc9Uc2bgFz
im6ly5U+m103cv+kJbTA7ljzLUj0sd3kDY2bWkGW9AMi5RBHRB8peOKfYB0kYW5Pa8M3FnpzYDuj
Jm7ve3DQGEALXLF+Rd0PtKLeTTLDqBABs1jRetCSZOaq9d4TbbtbbQWra8LxV+woVHB07OWwaV/5
pZYr7fBRJJfuhMzIrFtdeXuUv3n9i0CUJ6f/vQSzggR1/niVB2sOZfzsvG9rnpXtRRGMgftN46pC
miKWYfu4RIK9MzNCYGAMud7ZvXs0jXZEi8obI14eA2RLIBBXtCf4R1uVDBtGXAG5uxvJhTQfCEIK
CisvWFSbEMMXwiQ0AkgfxZ9txpqre8lIA6RQRT7bqsc/JydQP7qgqHAssUwNu9mymGrSKlCFAf35
Y5lcU19CBmaO1XjipF0Y7hFxZr/xmU09Js5hxc+C5QmsFpuYPNZBlkdj9smch5oRHqyMBZl4st/4
7VnMmqsUJcD0LE3Kxr5C39bKOxQrYePTcK0iFNGQV6iKPpL4e49jEHXtFBrKuLHWKlxNlO88s33R
tWaxwUsS3fC49/VX1F+/+WHiZHuygJIyBtY0l4EORCg3vqUiHyoYNJl0CI/uPh2R/WV8i/01kavF
1TRZQCk3G24ywyB9fuvzq1uRhnn2kP+01yHdmPLuR0sMmZbWDeUWqBa5lYcf2OcJhRC6Zx5+7O/U
AFtgkCryY4ZjAFbpAFHSZjMN/EoQjC05k/aJnpxShqvv/MpJlpPZpBWEB56gFCfLcWVHGRoq7+Sn
3wFklhR+3kNOBQCZePXhKbOEN3Xl/28RswsOp7dsOU+CKH6jfCuV6tk3e6LcbjsJI6GpwCdy2vvJ
yzaQnTYDy9nOedEZK7udNLqeiLhoZwTmMTJFKmc17BC3aAmcf8yuG6sNnNk52ZIJ4J7LdqEjGreL
VUSWBkAj9DEiqBEu+SCww+eq4MWcL0SOhnhPuFXCrnNPD0wJNu7CC2SFsO71B2AUFpv1NGu+J4Pj
cDvq79TaP41uWCV9UVXbkI5ElD2tUqKhc8RnagzloSXAzNywhdLbi+DHnxEsIy3a8uLp38upOAEY
uLqDHUURnzRoDRnS7dH4qFtbLJCqyQ20WLxxYwD5LEURqcAucApj0eRxZ+JA1l+4VLFCJWAffb86
Q+WemTv/fvYarR3MqYVj9WqYzQPX7swW7eyUS044dTSZIax8ke3wXPTcuO+OlOmo9SPztyDnAtXp
AGkp3vTBzwZ7kDOvQylpVAhov3ZNTCENrnlSY4Fty5Mv4NQzwWil9sDpNDCKOFv169+zR1sI3CAN
mlt5YW5kuzZw/dA5kTMZiMqpTnAawft7zGRHnKROPK7wqfV4EsS2eIkVUhrr+nliAGDl3NqUf2m9
hOUViRBLYyfGlQUoy7rXuRPk7jOcOG/c7FdtUR9H6x/sENcSsRio9Wh3DJPKlplCL3TlLRdqAhHa
V1Bh5xizhz9DeFRSe7SUTusR/GCHrvkBMuw5BD/RsV7FZLfqZmJhXUh3hcFhOuVwQDq3K9xnS6QB
NKZQ6iT0wTiGZRpUksHp6QadCoREfjdgheydd+DXhfL8PfuXrJllKxJc83fbnOoUBA4dxaoBKsgh
8Jc2plzKDxO7cP/oSewwJdW1HHL5xZRSnPH119rawHG1GshvRQDRXS/H5nKNEkmV32zxb58KKsx5
xwsyRiO2uaTWtYFJ0BZ62VhsCjozmjCIWU+ORZf0euslfIoLxtNkCjFI8wPQaVNj6wkDDpoB8sG8
eKy2eIUX1L3gNm/4fQoyB4osDjt4FS7TqKwFbRREZcvg0ybnziwyndXqbgyIO9XDummKZ8PXyMWq
oLX3zcWltgH7hB9MxTWk1un50Sz41BZodFOKmuYiZFSVaeJZRIgUzI+I+yPmwHZgRoIxfyAFxr7y
UHkeaxyZ3YE1MAfZmpLF30xDcAvUUmZYVcAtwtEvCFLqmB6UNsR2HGrxO3+Ukm3EIIqGX8P3UghG
qeuarHnyYnvdVHXp5PM+GU+OdUmsX3D4cy72doPBy5TZMRAOAm4l7LDO6Ry/mq2BCPcYvZTQ3kiL
fh+F6O71k/yCBfolkD4UNcZjqQAqYjL3PAseQ1A5NqdvhfGhOfBTATO7rRIBVcGBs1XGpBNf05Og
/EBUHrYDKRv0HRLH1oXePg82zdkunyJC6T5pCzEYstbJjGbAQmEeDMG7UJGmRtq7bNvLFVoRyEk6
LHriA5FwPLPa76rMQIGDm/7y6a/gWWz+cHWSTGAJ+bO5TOUmJn67AnD8IzuXdtTAc2oH+jBVv/Xo
LUgmLAlySZiWELbjJzngLFfPMCvHdXz7XbDWzXYPYXn50XNd/JVg5zSz4tKglxe0bz6MtARGuk+q
AzPBRm/0+LoKTnR0Y8Lo0gNr8EE3aWn1MqwIj1tL99OkbtqCe6bQDYesaFAqIMV/Cjd0Yr4zgVhN
rCNnHsVmr1Bn5iOtIygfWX0UNb2BIa3uT/IiWR2IabVRr90dR/35TsviBMTRDYTWjamhaLjQPyfN
54Su7wQMbwg/3AHjKk6UcX/6Q4xrbFr/9iombD7Jis7XHFdl/CrFu/T7U3RHuUmd/xzTEu0yurrY
mN9sGn74p8nLhXYoNaNJQ6M+xeH03zkUfqozSHVmdnh8mpoVkplP1TqIPOSqWpjpsE+ZyThCGI+0
fKK8F+2sZz/pHdtofyzZH0u2aHbhhwkHR7pNMXNM2wuJ5AoQB+k7ZEFnh27zmqXY7FLdGU26CWNN
hz7EcXM64Fn6tLA2sQVsNnUuvBOK0DkM3virlNUy6FBla8EN8XJYDZ6o7kPMlb1llVgKvfDxAKzc
ZcBvFQ6R2wbYGO0qFRYQcPiNeGxkuU3ErWVPdkvRRap1Ctcmc8CCiokb/T7yiJDkr6iMekr0Wg9V
e7aZ/KXOCcb8lEbc9UZDqP/BACqrz5s7/HUuevXa9XAJlOKLg4NECQivh3RG8Oapc5NFMlw1wY5O
vW9WGkjlP6fvVw0E6FYmcWATRBueewng4dZpwr1mT/5qmqnGsRLQrLWjZw5JxfsCjA0o3nlBTUSK
Tc7pyzc0AiqPh45lO85KEZegjxJNQ4eIVgI0qDvxymnLUa1HZhzlGuReUGUbqjSAKfQhXvPDo8b3
CK6p9edkRr1IjHHfuEfWodyy+1PElXgXPzql9UQX1aBnugLy9NNZOdCooqpdMnlkrd6bGJRhpmCc
iPBN3y0ieGPwgZ5UM/kmXWRfuArMoXvlepYBLMq//sXtlSCJ4QQobYUkJk2A4VnE5JInpp1+pAs+
L94un7NJkD0b0o0viRdDFOk2UlOrBmS0cwqNcZwhEK1uL4J7dsBSBT5FEX0NpqSjs3dkrz1KkhfI
wmYPsBoqeVEYdQSV3j+EjoCUMo8PZ9w6s3BexFJTLd19ZbznkVtDjiHKggyI3/L8bvhF2bBQvbag
7oqnZpq9UTeYNVEad02Mie7aA7HNMBJTUPzFvVjHXy1Ii+a/3VHnJQa9jsC5MI0u7jKhM+Ljevc5
PoYkIUPsm0aQqN8jqCGSs6F1I4hcUoJtb0V/sB1tTmx/qrBFrYEC/1Fl2Vuofb/SQX9ltUAE0DxQ
H8fnSOsFvJXU7SAGJ7MR5E2fqLsMD99sJYPC3a2/NfEKgXcGUOoVVp9Y2FsBiVNBSLRxSPNu9k5O
gON969SrcssGPdfxS3DO8xJU6+u/Lj3kgg8vl7jxit0vzEPyJsR+O9CTqL8DWiGsGug9McW2Cam+
xwKFlaisWpZqUdpL6pJJVfxxH+TkodKPY42ZFTUD+YgMIZwADR9NyjchlyPcYNakSKqU43cWqirV
Qr6pTzSfZZ+ZYf18sCXHUN2yzpFCQQX6b+877GBTw6NAHIafR21JJ9O22iYHcUgKRobl/8a8ecBV
kIaHP6bB0D4cV3V+0Udfdf5wKzrWlBLCbkwolAc6GpNTK/lXCAaRxTjpCKObadxEf9NTHfWQAZR3
6ktyBdf0gi1EgeIpxvvO5SQ8bqk0f+bEcLKGqKDfeXm63Tmr+gHT2e+4mTJeCy5+9rlu8htFZMdc
fGILCLkvSPJK6IakFA30NkGCILhkWWcn9B7cWif2nYZDyH9nUFLYtTvWIOv+wBR5pqIsiUf7UMGs
9YBySHp2lJgNnCjgWom+voz5SgT0jDT7EMt8pI6AR25PmVT0C5GSfSya5i3jdibwBTi/z3JTX+9f
JFeY73eokIdT2AdNPK1i4Ihum8LHGuIlEPrK6+/mzV1FRVUDGz3f3I2xhK93op67JWpm2nXu/CdC
ZblOJUdiZhs5IghFGL527wIhdAqghJYXJIscB3etI+ZCeNS/7IBzL795sFp+uurNFECTPcXDaFws
oLCulJuRhHHRFIzfKZKSMzwGk4yKVD05T3eO+ki6ejOQeYfbm1SQt6wGZQ682KQZ9vWf/AJJAEQa
4az3YkPRRrl3S1/nhzjMmLZWPyl522oeMaQWHAYXPessk0/RxB9d7mLG5TxUBPogctn/ZtwicaOl
ryNe6iB1O3giJDO+slab1g1umYWxqfW4H+EJo/2qvgkY8BBZoDB5AWley/re1zYbTqpOFWJaZdLj
EbYqeG9dsp8cNOaewGEe3wrvohCkLv2S4gsUp34O1K98QaHdZuaLOGt9xesx/EgtR/DL1HdZeoXi
Ioh61tK6De+ZB5R9iiI6l8VS1HjNFxK0vPPh5/Xyi+BgWlocBf1bMSpZBRIUl48u21xDDjTqKesI
zb9FsBnyYpowmxaENcRlqwJCoMNC/X4yXrLxK2fREiLSe38OpCvh6n9YMakV6sy988LZF2OQwgzc
mkVWiguAsl3ksV6DDVu3ReptD4bDtETEAT9U3h4UB6dW1FpfHYf6KFF+XWtRbykQnfIEFAtb1SOt
7w3AaT0ghJM4v8Dvljdqc5JAhTSc6aUyVGa+kYApT8/sEkqvNmwSlVDuk0pMMw1HnfHD+AuZoSTu
D8R5gMwmA1VGQymXqo2CVXuLmzHFktyD8FEbQnrZ56tEvzjpf6eqF8Uy5cT9vObe3IRGpxENf6W5
dsGC8LcZ2DbuTtPL+t/l56S+/K5Kx/ylkTFMpntHUny/WfTh5kV/lcnBu/iKYcIJVcfnP7NYigxH
RohlMgKOOK9Te+V2HNVqrOPObg+gRyLgRt7s2Vt+hH4LXID6Zy8Frzz1ujSA+CZ7wPD+02sVsCGM
KUdHSt+bhck3r+uMNe844XaUOvk0uFLl1heDSif9dnb5WUaAHgLSAi9y9iljU7k9RWY8IH7UoJsh
47QZQMfQzF7wD1Zk8oGtHAD2h378VA4ReTcOxJWjKm3L9JNBZsm+dJ+80AMAWawlr35yZJpIrjGv
Yf4VNLi9VT4J2vE/X3iHtIJXtH3nW+oGQPX77FRXofmaQediZkzirlkEXFQvbHnApJaZwKXfW1cy
W6h97uLnY5yfaauhSASKFmU1MmuwsUyeOtOg3GTCuqh+R42g1e5Ap2LdKKYXb9xupGvSwEnATXaE
0i+HWSPgXaqwHUM4auCcDSk+kWvr6h1iZcxecNDakHWYX34OTYOS1BD1S+ll9dYeJNmuLiCb1lOz
D5d2vT7k4qJCbYAn2rU9GzEG7sWKKCgZu2Yf8fbFH7l1OEx7UJ9TppZizwCyb2Na6ATDa9wQv21X
bNN0+SOtKNGDaiPZxYIPUXqFR5A7EQqEv74gcM9tRzjpvz2mWxhB8BrmCoq+AS+dREQi5ba3GXHx
aptdQxbV95yua4yr2CD7aBLDqaRd3jFiNWC/uwAYQO/Av6D55on7GV1XV+uGXiwsrZpSbLsOCbKQ
kp4uFiYV/hNjY8X2aRIL8qcMKBJkw0hfjBCiZTBwdKdWjRaFXTYJfptSpukTHhuxlGPRXIcEYb0R
nTB417/3yQBgPGsbX5AlValL0hvo5VxCwitmjZbf+/bbAdy6FhltHe66d02zBT2SlXJkq2wmVP3s
qJm1qIUEQNe4x1NUgepvynZuR47mm2y7S6U2MTDjtPhcUmW9VQdea+95Lt6pU6xum7w0PkDM1dne
zjIkMzLeODm3hZkkeE1NxxplJCE/uxf0Pz02DE0tc1+1EW61Sw7GioZa2yyV1+gLRmKul3VOcQ7S
7DmNnY4NHVgkthgKWdlzDzKrd3lLvfwv7GTwUrxusMVgnc1vCvb7o2P0B3bl3CvzwNCo81Ixovta
IVq9Re+wrLFXQI4di1UBheNBVvrAaER59K5iuJESf9RVQe74PaGVzkLetFGwtRoUTa0zFK/0bg/j
JB66P1LLWhMjQCn8m1p/0CYWlPIIShPOqWWTdrQ1mqvVCfUOhN7MTo4FXENagDRg1geeYHzg9sm1
Yg9qu0vpNhgEjJi6l71qBePrAnXp0uyyh4cJzj0UOCIGKK5BC8uIz/TvX1qa4kqYlBSTQs2UZPAf
ojvcFfGRH4AszO0/YC7lGAWW4ILBc2DE1FNdZgIZeDS81/uNpNCCs92tIy6KioaeabJ7ymYCCHKe
6wjbGWggSZprlnnCMfop45L//7fEa2BSs7rOFFX64YEgoht5JcZXyloSuebEo9ZRpWPRJmNP5gti
6OfR3rnMng6SaW6gsDUwNt2qWpPbfR2Fx1AQlagvaKMRn0o3N0U/JVQz5wDPk9dfPMwSI4+oaj7w
7vRNjPBSmCQ7B1+ejCzv9Ty2B9HL6lc+bCq0UJv2BuF6r6Rhvv5CReTNro6Dt7PdNcnp1cCRB+aJ
c+Za9TCuen4Fi8W6xvSajDbCoc0WpK8cpU72GIOnvja1s+S0cg9H49u7ld+fTncSOGIUJGkFsxoA
x1yviByTPmDp3MmGtl4PdKtOtYwu1IYsawJz00gG7a1FvZllhT/s24TvvMKUgkgAZDfSCCdLlH7k
mjA7bgNfJbuRclyJ6PET7vwcJeLGXVCFnbeLHYTcS4tiD13XEVB3xOszJJo0z8mRPo22i8odWU36
RuW8OTSrz8ylkTQmBLYBNPgEJkTM4wPym/tLw6TbZ4pF9cWoedVF1aTiLQ9HRGDUqVy5VIiQsm/8
2A/G0CG4D0zXrsFMwy5i04fkt2bAbyo71m58S9Pj/Whop/39CxtyLvncCfo2rPSenF5nisDn44Os
OTd6ioVz1QgWgRtH/DkmpLdRAYx4yn5H9xRajgDITpr3LkTbRH1VTZd2vHtjgSYnUQ77kxlN7B5P
/mdm15Oo1BGNFPtPy7RWKQ24mFSLZnwcbI2Zb6W3vJv5gytzw1HgQd/+p4z64BDYXuwE6o4GrGNg
rRa79+9DcfN5T8ieHkZa1bNLk3qr3qbjUj36wjGCXGTaS59Ld09jty+wjemSpDOHwAzonoMxBhuj
X3c+oKCgQ30/Dkc3xF2gQCZd9aKUH6GjNDphHXL4+Hevi2OuelBuBjztYFHn4Nm0eXlqYuPsDpOV
6WBPPKs/JrXcTcIE2kOXfhdoUdSNjRLKk4OvkYHk95ASfkaXtQ5QM2iGmAMFxkZ71MY0ROTQJfbg
elYedPkYBN4Lks/JG/BphaesRBzvExCB8Op3O4nDnJe/zIpM3pTnHIyng89EufNLdBeOS+UlsloP
Fi0XuzWUyxRrV02ADkyZ8ldlb+j2yWTZsYgQ9a9oZTe1MzEanC99SkUwlTXxGYne80zwlRuCeoCa
XqoPmeYRFpY3vczIz1HxTPQLTKwttUzpzEBoGJBROJ3PimYe6qbNOJ3ZZVneLMZ3wGIqfwIrj0HV
7evGxqWzccGPiYKlLwCCyvMMmWTp2oZeLkeeS52GVevKpCYVsb/4h+4PAHCT/v3fWoOqWmqwQgL/
xx9cAs3a/9mpU+ndJp9YxDJ/tPgkJzjbGjHOOgquFv84HoscfUiaoyrEaavaNUDHSUVBV1kkSQnR
REQZUbTzX9Tr0vDlf4lNT6KgBV2KlMCXuCaBvl6Tg0Pq+jZoid1OJ5JIZMvT34hiRvt9cb1oQRbG
p5SkqD1sWhyOkwX59WvOvS5jJMgQw/LsCp6peVWt/NWUjk75rJIzvBCdV5BK79v6OpjuU0HEAKoe
AhNNZrbVddyFbxyUzjOXBbnClN+91twC7HCaVyid6vnXrbDD0n8DZkMJydtQD3JKNDfQzmVWrmHU
GPYQRKGtLWOx20wtnkSiBlZbyUHq91se5kAVadvUkNi3rpQZ01FOZNb0J3LTXC/0rqPN/N8m5IEi
yEJc/7p8YdZrmtgpax3ZIR9SEJFlq9x7H/gRQH6IMQx3zzkwQaCiw/etKokEzgii/cZi6OH9d8Pu
557MDSejam2+sTozcRflRROycf50nAwZkjbwt0ImCCo/855r4AWWVhG7HKzrf9ZCp71b8kt5pnjT
uKRXyc4aDiFykbjerRvJsVRMqy6Gxke8W8EwKy03VMNPWWU+aQLrVVarAJ7NrdpBusefanMocCNc
ykeERH6t+VtEJJs/D3TyYbklqA57ZUMAMXgUuW1R65O7nwvc6/CW7pd54NINfR6mASzhT4QIMkhF
iBSHW69a+x6nwlkBWJkDSKWXpQOKpv9vnWaC4FHJ5rs3Drz5iekIpummI9lxXmgaIvLErd7Cie79
cSImmKJ2PC5iLTkEMPphfqYSedKyF14pSmVcXcc56LjRD3Nc0ABEaqlH1eTtcjUEG/5HzhFME++I
uHxTCqqp3v/4fHvPH2+WNPF7qgfe93VDMzthJa7r+3Rlv8jB6o86owkLyq93XgfKDtKzPpTyvb/d
RYxZKIJWPEBudJBLXmNQII7BO/g5RY7WRFHrE/z2ikli4Ti1/6GQntxrtCN4YdTWLv6OPHXuBDiO
UmeNU/mZ1AeLrc4R3xzrecedkq/sFVB+p2lAYwEmwhmuKvV3401io0nSlQkQf8Np9iaUn1gYc+OX
exyw7Dv40PPFWTMENBRnapwpZgbDo/cao/1J5bKuP/z5hlDd4nfTpwuP2RQlhVVqOm2J9mLGNoir
tbkOai+qPtwUbGlToCo7mLpFWApjCibmzcJ2f3itoR1zS/99Oi06ni4Akx6Bf9KWPjFw/Vioan9j
p+C18HXG0nn3NNZag13guMh+kDk/3JdMS06+tbM2OgPM3vxXXghctXnBv7xzgd5VG18rrwh2Datq
GznBP0xxQJPQnVYPeJTG48XCge1zDbHWIPzLe+BWsn5weXdVQsVhQtFXVWZWXldRsShxiEriI/UI
JpYzhF/KXS34YEknqgDVGYFRF10YUPl4HlshBQ0fC6PA7T37DvHW7SNfvZoMU0EhMurxr5Qxeouq
wjwwtvkRZmOFM21lwNXIW5iNw2YUIFm/PPBBSLo48U/2CrZOIMgK86Ayx7/ztIIOfnFlX4oVR9X1
sFk1rXYXixXEk1WL9NSeQHGAPVfGv2mvJiOIwT7Tmv0a6SL6VnTf7EQput/F0EohbfGaYzyiX0wR
wvgUsE3N2hhwvU55nEXKWHhh+nMiKCuqkuaBYz7lEWGFhTHi8qW5WgmTlKzeXfCxp+AjSpOYgVtm
Mu8Htdv9RGoi+he69Tgw0B9JlyOU1Vv/FdjupBshWWpEOIkcFFWAMmqLKWU9pv31FOeigoMlppdd
8bbkrkPJhWVFIAsNewveHH9Q3vbmmkv2PKs3I5shymAFjaJ8mYlY4CK4kWvu6kmBkBxpH0td+UUB
9LPzUPvv+OgJlx+UDUiUNDKG2N43V8g8x24wHpKd65/F2/YMXm6BO8zLMlfwOBPEx18dgI0WhOXI
bNfywrY8BqKQDxj7nGlItqAx9XpbWAqmRdGmzwU/UbJgf0q+3LOW+tlfOgolO1BS4DYWhHMzyNVw
44hNBJYD39rcL+5jW+vlaEKj2R4zQJlx2qrgTkzu3t9nr2yrqPL4NWkVfRWEjNf9xNy2xr0RmClI
dTD6EGA0qMzU/o3k7xt9DGokHJt7g0I0pZft4fWvL27KWrZaxGyzEQZMfEiHtgmicwbkn2269F9n
e2R2IHQCoHz85xqsvO6gVO2lZ6/CTpl4jTcAhUEVVEc5kG3fH8xNfA+pIowIpUf79hSCvWj/GJpp
ZPwdswm3s1gChQ2fwDC1vEMiBnzftG2cWJacvQKx8pyyQrYb8umpJYTPfPpyIUog/wwPinDvy+gK
6sYt6AodIoFNL/rEVS6a+xiELjlTBxLpikA59gmZ4OxJubk91th6OlZzQPb0QBKuddQ5lvhFT1er
OBEyjkDUDnEmHLRdmho8zT7QEguWZH/ls/eLnq15uivT3XoDNo3Ti2BE2faETOB1ceaINZg8RKTV
CeTwZnsNW5kGJHTUUvn0cSa6B6JEGvylRwseC8765DjRtrSHWNIACvsHNxnvvCPXGXyVdHIlkTKz
KpR8P9sysjEfwl4oKgLnDKIaXRER5tNxJM6vBC0OYEZX0f6Vgc7kSOOnXv1/bckWruZWwDIQggCA
qqUwksMsCFCyBmVZ1okEf9aGzitNF7VR3A+J3qNGEvsM3WYjKrzcEXaeiwJStSTfP0Z2VzCfF2Zf
m2II8h/ryK56FFJD+YLWRSR2NxotR3kQZgAbfep8KRtWhvJW14IksIZHAC1C84Uqunw+01RpcZdy
bfdy6REEUfJYhhZAtjT5lk0CSkyYYQwzvE/NypmGLB3eR22KbgpUs5G3vh8hTD1+2OTu+wqsrERl
yDQPYiDIq8oYnIKKR84BP1WoqT0EjaCLxND1wjDxwQvxkEcBnnMOi0odN0NVUrA4jzPPs6BvbnHS
igBlStVe7RRTF5I+Hn6aUsNSrUuKrU6v6hkG0gxnKxShxuMS5fKec5rH8eePq6RhJ8Hkdo2dOzUm
nVc6bjZSaxb+MNX4B7N3fpWhqkGoM1xxYtRLOz4x4A66iZsS2hSLBPqwOuKniHKIL87OaccWlU1y
XKvWgh0L4n+UGwDhsTo5pPwFrdtIMSN7rkA42vxO+FIOBjFtNjWT8aNdhwr/0ESKMSBjbttTWVMd
RXHxE2g6k6aah57UAlQmkEVshkaXdFwD+h2Dwrai5FkNTyJV1l7iLnSZyHN/NUWKuYb/MBBP8nha
E5lhivpRiGkePxrwrMAeeSw2Ut70MJuNfPWPQ9jXAHf9gHFTj22Ll4FQagi3NsU/r0wxYKcjTW7t
5nFCqgrJmdmJaDfkcv0w3Pcwm457yhWEKplGBCVmrIlmw5ZmdiZxorBBPMTaUajBArtDvQwAUXXr
znb1Q/Rfy0X43fXOHXpVlckjdFROQ+iCEwCFPWG+EqjhrVm0d+TuhLpi8Vq4LgLvcmNwQzhCCF7B
PM/JhiKrDv0qVgxmdnR8ju+72HW6/NuCGRXxX39kWsJBCetcOtdrEGYFsGytpfEwPl5IHy6hFRFA
HobO5ZfZ9BDzSUi1qtPRSOTgC9X6HT2Q0zmv8vjDOUxREAZSnLtpuas/RbJl2a7cYmrEkaM+BBLd
Iy1OdXgv2dbHygH7p50G6xxv+LJriwaHpOXb+cmQF3HGkvpmFu9VU+fcAzt9YFkk/2SwO2B/JbMq
OmENIBt9sJEOjHsOIUL49f/5by2gpF3EVToEFDN1Te+48MnQtFIU/xGjO+AeE/q9wyg2at7mPx4c
pd8nT9Qn9ruwnmkZiMTaVmorEmodbRmJR/sHbPqbikPRyjt11OgV68rlUjVVygvRbRYxMqIuMAlU
D7JlrkTRu/YnXfsftsd4nwWjNWU04yRREWLfs/RVFKu7LA0vUpLr9QM8pUJxWbLYZBp4rPHxeZ4l
tWNuyYhlt3njg1qFWhHeb0OaQJwqP9jl9V/0MuMkKYfvtTylvVs8fS/hlQ+eham4RmB9oO8redRm
vvbiMCXyYXc5kS6DQorWwxKHwjPsNfw370jXLHAPbkrl+jtVqqzucydPsiAAVrCIH4+A7m4g+CKK
jgZVDdfyoVxg3OEs8RSbQwqXC2pRv/s3dS5DDVUXDh9pOHZ/V4N08LmT7BJpL6JYd6dcTQhuQQvI
DS030BUzicR6hWTWL1JQEkfseqZAZcIh+cKLhHcRkWu/4Qu5oKjfQP6ovC9G+WJtWy1he1XT0GZU
Tbeysca3ehW6EQ1A294xHTzbUf144RTsugD8lryvVRAZhEkO/3pY83nyIJW0fPyjT4FcPHH32E3V
HLg+7udyqaVLkzYqUY9QIQxa+W49frpL9rAlD88Ypz/e7Z9kf4Z0in/VgrE3wCG8vVUENqr0zXXN
jTT8qLQk6sqbKdg71evr+LpCCRs/C84EYSYgPQn1PJJMvmYbvu2cn2d1mMLyWs38O+wU/d6ONfy6
xPb+DSnn/mD+lsFZR7tUxC9sgZL6xIfS+RPsombwp2AVVfxx71Z246AVZZ41NZK2NgciuCJuUT/M
QXRNRIhz7JxXaYWmALCLPQ4lJUWyWzuqRdd9DKNaJn5xJkCNmc0sQ1ndHAGdzXMRE3pLwxFaqlA5
e17GvitQEdkCMBLBUAQPU/r6YW6Q2q0pYYgld1gm2KjQ1K7G7PK75pL47Bdpnnm9j+DEP0X/NpJ5
bW05BFM0eH6WXZQOIbhgBndYDJWVgqjGhafZlbgZFzTPAq8jO1AkO1B/O0NzTGKHfObyU3Qzf8k5
1qWa9KCR1CkY9jcreCsfSy00nouvJdojmHjQLU/jfDTaTAP4h7T6gkYB7oNl2Q/diHn8Y+nhImWU
371MRRjVxB7Ax21ilMMAEfEQ2tyUiHyMS7an3nIX1ilZvnOjeR9UN9oZi12z1QNVvPEompO7myuS
3l5AbCygCjgi5nJSpaAgo4oibNR7TmdX/Yd/CB49FwUcbBiKu1QWmjnmwsdXPvOHAD7/edhDUb/v
TWN8yj4J1TzNKuBCjyCUKWiPOb7Y9ivAMDxlSLIZyqMiWQGwhfeBn2nbWjJPbFCeubd8tQgKxXCF
/azIrk1nMwIet1dLohtJ091ZGK8JINE3iKeqsVQIuBl67nCj7lz+X59Ix7dgrTvQlP9z+lPSlUep
BDzVsJf+lsljYXxV3kHMdG+UyTEQyXhbhpT4+nlWSi9WDkaRb8fzei8fV5XkzdKdQn0mayuwhNq2
X05gJRAWxw38ZW9DDoD49HashopGsTaGn1/NVY5Uv9Jr/7FWxHryrnP3/dg4W3UAt+P50bOPU+9z
5L+oQMvKdut63ARv86vNvthmd84ntiBi397tfCNNL9KVNWJW81i7TXoIn1qrvJBE77701aq+EErY
9VgDDaf+mHHvH0YAm1EFjoffuiOfP72O6jt7eRvAgU+cO5wFc87dhf2zA/snH+ASw/CfYEkQDv0I
b6OL34k5Jp1uJgLUXYNQeq+WounR487Kj9h8qLydDpajWWRDxL+g7gIUY4/lL/TAcIuSG+3S6u3q
o0ZoRe2SAZuCSEma/UqCkfKlnS91lDOGUgIJCFTYq8XY8lpjKjE/qJF/QyF/hy/ApGX5nRPqfELc
plCN4RnBXPRbuaL8+0joD75aPjs4cmRxT9B8SZvx42xNZt4u+W/hyj/ORX/jG0FtG1Mi/hORN1mD
4VSV87a4ErFQ0K5CMgoevNox3XPA+ZhTr48yFKcFOVmVXHQq6Lm41N0VoqvuddtLd80aYbE8hByT
6bLUrYIgyiPiMG88X+XTyCGLv5ANmk5dna4zRVQnjeDSTCm8d+Y+HjPQ978Vxfvvz3IsWRL7+6uh
MRcRp4cRqFMqUlhwXwSXMupsKirKT+Z+H0raU+PDOoM9i8Li6yEJ3aF1ntlWDOCYbqNnUk+lVOhg
1URfvJMWuZlPlDAbLoRBVX7Fq0ZLyzZ7k4veHXoZMzYTlUhv8cLDgNAZqSAgHC7NSqSGN1FwrQJS
pOnK8kJWYa3MfVuTJD5I2LQXA2a0saRHEsIDoAvHaJx9Hme7XDml7MDTj3AxfOLeK2Z3BSVE6RED
ZFvido25YZD7ZSx3GSjsiIpDgKp+GSIRzDDXc3HYH6vSBigpmSdq/plQnVXCwOW8CQci258gPeMl
GJXx/DrG4//aQd1noLNz2ECms4yaRbI+vqv0HqPqPL8b0X3HxYUnUsqnd8CGyAe1bMPwSVTNlVlw
YFY5ZIK7PQ2gcBk0SuPo3oOGxp0332yvSk3flYOioa5FR2nYKd9cyYAFAjD/2tn1vRRy+bg5OWKQ
0J8NO+lIO8TYseFeOWh3uIMkcdUEmNHKKqk/MdJI1xrCw3p3D6aznIWYzvWd4mIY6QbJvUEN9fnk
M/YfFiDi/gfDcdglPpUlnwwBjGJIY2Q1LWSBVGLLB49+1FQ5fUWOjFQnjGNabWV09suRNFrDfofv
zVcorK+U7j46qb0DWcfuSDJt+pg5TyMF0H/8h9y4CMfxWLxDQmu6vfeR8nBFDIeNLj79A8US7iLl
efP8Ks5S+qjD55pzyFk+xtpdziXsfNJFxuvdqc+Tvpo54T7Ac5SoQUkfmCVmhQU9fnpIciTuA+LV
nOjJ01undSDb61jVvDbQ52xwdR+w27o5Bd9QjND6+rlwJ4zQu2I8QCDl660FAKlPt6WIO34c6RcG
j5V02DS6aYqsA/sYnafpKmaEFXR8iozqF++iRvuVzN5CZ8ySn1mL5A+kXOojuYLgLkGQAZ/aX/iI
IgBB+dsxfDK9lynSb8//q8Zlzrs/ZFr6T+F49o5RtqLBQTclBFkMshPGyGT9XO5kr4WjyEDWNKHr
/Ryg3D0A+pzhjlj6H+IxqM3Isd7U6+29qkhRutODBWo9Dwsl5GXGRsHdAzHq3fUXGBQ49Qf5UR5r
hLSl86hDWItFmWXvzjbLt44fqCUCWILr1k5XqwnW4EnVDSI1XaJD6DvXKme1VmauGwZvBRvAn12t
s0dGStMZ+c33IxEIvdUbvDJHuS/ax+LSjTEG+RnTYTyWv+3LnyDVKnzbS1cRfabApZETP3c0YgeB
EindWzAVLSmrupjkApuEy/eldp49cmf9umQRQSQctd4sQaZAVcdjBFl/zBZ1woR1VtQeqzKQhao0
tyF5IFrABLr/skmreQMWxjYacY7dmsV1rZnZJC+lPy69WnPj0mBGIBPZVxVJ5S2DSW8M52V4WneV
UFNGqBndrWZymZj9OOLaBMUFnXmAVz3QjnXH9RBcgbT3V0MPtFfve5pyYKixxtrwC5Sk+Df3mRnT
wEr0eV82NFJI7GXaSnYfshlBZkZ4nww9VgsMpmomvfDlPYTwAQK0xJGWKyruwlg1WLOPjynY1jt4
aIr8EwV/Ab2EkBGrPlYM9qBS6TSR+YRPFOTT312ksZBm6QE+oq3GqAXLGHGEb/nTtW3uSaxfAyZu
PUs9Z9YlXuNvLye2EnUsC+/I7bcslhukXcs/DlM/kVNZXC/MS3vlWYYMwozNn6x0LBLtwzODdn7Q
MQnbVnjhfxHXRezlekdg7HnlzWi1hh5tOBqy1Qr+mhGeM2YrRhQd90DiARVcgtq1vu7LI04rblKH
krMjoF+pCo6klAOYgdq6hQ6vTwHKoVSYcpS48dqBFlr87dSaovUGkkIxyNtCgJhOKq2HPN14CuNS
lxvSN++2S2DQPz5uh1zVjckBxNGPa5lTiPCEPE/DP7xhQYTOBieR85JKdv2VvAank6K30FQpNixA
8N4W+eAg6UWLjLdXrkKNVDmsWhzrfSin0pdeze0Ko4cpLu8rR7hDnDowF3XgjEfiqAD9s7xJcbmI
jwmzJrw2EbnAJXqvfbIW7JcfiNLWR/zJKqS++oBTjwyie3AFBiTTX33IFD+ntzfv12B7nRuegJRy
SvCCbPIFRjOHSE1MtenJKA2N8lr2HEv2DAdvchbYvcNLfsgAlbTD0UM/QNZBbP6j0mcUGoeHerr9
hi/QijVXqubcuUf36LKZ7Wo1mhtQvFcA7FkoG+Pnne9ocl2dzhpZMDJtqU6jPQZBgFjwpgsrq/Db
EeZ+Xn+iJovxZD/3IgVAtt5JXP0hjL8eZGyc+Muu9gXQGAGDE2R2yCEO0/dGJxdbq+XuKtNbMmR5
82abMMktMUNpbrT1YrvRW8JULGoXzYjCfMXON9A26ryyJtTMPjRvJMDIXnHmQw/KuUu96tXdw6P/
PA9D//I/Hi8esrR9d35SEI+UrdlZLcT8WVztBFAQ9BAGPc5JABUJQXchvOWpvaz9y6y8iijunV2T
C7VGu6u1atgRAKswUtMCo9x+twyZWbAFPkFeJhj74ThsRD6TJgt5zhOWT+7l2YAhfF5t17QBIbYE
DQ558DMHJK8LuiWIULzWWAA6rN8jTHF9tV3ucOgTjoE9JRe+N5+gUVxKLSBObtl0pEgL4sW3YR1z
l8v67EDGGZYcEOY9WzMyBmulUf3XVVa0kkl9mU3CltoJABkAgBjbIxKxnt14AnQBw5sVGJCJ52g9
ger2qt8WmPzKAIVZA6TtpkLjRZlnvhiLsLGkHabcOtEMr60kLjXjBFKl5cNlAQb7iEKBHoSeU8S4
upABlGjlB4HwLOdM6ZnzibVyu8Jj3gBswsrMNmL9J5z0/ebsez0nseTkGbCGp1r9n/Netrd1TSsI
OTMtHTeP6dN7uhjeQTcgqOeE2lN9nHyk8r4zNFcgI/oeA4C2xG7tuVhtLmtU3qdb7AMalalAkeNG
0G9YYmGxUiTagnD7gyLK3hpzrhj1wSRj8DF3NqDKrwiwMOiCYgyrWBNRxssq0TVjmikTn9tysYQm
3oH5KZ1CdKMT1vMs37T1tRg+KFXf8KcI2gq2KxFmGQcSdzj6axV+Nm3AeE9BlC+d92P18XJK6DLZ
OrXbxqg1ykCu92No+6ZE5CC9MTLeRWFFCE701gQgN+KisNlQ738lFJUsOB2V9Jq8BrvkWA3srkb3
8SirfXphRcGB7KrernaRQrU+RR0gAyXrRSxW4ZLhTRL2i3MLNYx4+GFGOUp+30jHaDWq892hm1pi
Yh637ET+E+mgikX0bk1Q1vlcax9nQSRvQBJZgySvTSFja7iZ5EWO8qhdk0nvr8sVDb37M4ahe8pe
/buDXHlkIW7BtZiGDIolKZzEBpmgh1PrEvb8wwt+b3Ctnr3gH9IbXBug4Ao6yufyW3XQFwsjtj8H
av8EW5ftOsjqSBoAGnUS6XNc709z6S0cjEkxLQ2YSWY2n+QRiqeFXB47ZDnKGcTf5QPo4u/NyLni
/5Onl5m2gP2UzIcs5FQZivY4BdiGlxgES8ev1Y0EUWrp04829EfLF5D2qFOj1SoH9Ky8jwnzHia7
VbEuY8d+S1VkuPx5m+goQT4dSWGLNFTEXwTNKEm9adJ/PYR05ecyX7H8SzRLG4J7nEYADeAMPXvk
fRksUhF31pe6yS/WBVlYw/JVXUoxAz5Rmo0PBUyJ9CEUajVicfuTMOQmpsi7MhZJLQqJu0WDB7SD
PcJcpOrBEEwt5HqFnURFtndnG5Kf4JULRynx8pZoVI53k2dCxvHqGo5MoZmy1eHmdGYs9LJQCtjr
tiKmMaMNIFKzFLoqHZPN5d/2yPsELvQ9vi+c5x9//I7eS0yP5k/rHHfeGdMYuOiaDMDoQ7v+4r37
Ng6Dj8Pc9I1Fc6/0p9CLn0ESMcXg6zlcZRqEZpXzTcTk5ZMRRzupa/suTXQaGDDe/iJSICLgT2rh
VWicvTRgqN7iOFS3TlgL4YbhHNNfL/Tj6ZoJPnq95vbUqcJlDWVp6bnbRKMNC20byqKaHtC3zFU6
ys2W6xl3MFpcQzIru8qGw6J7tc1RRpXv1m395XbAFuRHykDxOiczlJfv4HCsh/hWWi4VBBoILorx
ORKMbhIxB9Zxr2JWs30OZrObiNrh7EYvnY1lKW2eZ+tjK5dC7uU9OkSyPtjCoe+WjVv5Wa1elRgA
gpYDhd8cYWGxrNLcmgi6mXuS0M5xFO1Bb4iWT3BwIOkRwz0HDlonIRaM20ddh2OwCt/G2WWBFM58
VD17XWhmweOozBjvVRtz6RTgvpHoq1mUSo4KbNqBOdTmxJb3mVEpw4FvVEPfuPG+BwELQafBXwRb
hg7DhvBVz0TEh/ie+Fs7zIAEIe44/c6VoHShhus0UGWq2UM0+ovFU9sa0+MLpUsdNHxmyoEv232X
1ESj9tvgupjnN1Yhbri2xaykEGHi+pwClz4RlhfVwKD4iXrh2/PcvzmJON7THtLBPywhMLoae9jq
hPvlIY/snaG+LEPt1Rp2hvijkj+yYA901HlvQdar5XO/NwYy+wHBnq83LpbzxdxPQgxDwb744jQr
MjZ0lepLIiFNNc1F3Aoe2DcAxGQUQ+QmW0LOtP00oVQPNWLlls7MUc/gLznNzBtCcl5YkNaDrCgT
225GBw1M8AOQHZcQMM/wVsO0pQnrpb8jKHWnf+R5O5povDVLpFFGaV6za+sc7/nq800/Dqbj/4vI
PwrlKszusiTIjqpzr40uIPuH17j/Yg5Dy5nFXsE4ZIyVd8t/192hkkEb8WDZZkilD79js9c43dq9
my6wAr24Ous9cnzVdXBiGfxVch9STVxHjjaBhMhSqPTMMp4hN++esiMSDjBURdtBQBMPPJRjhdfn
WEJ5Th6gEfURTLsGuxdIWPaiizoC+WeFRvmXtENf21NcEaadPlFxh6beOV6b6b0BLQ1wkfKHYBzd
EYPYiNcZ5q8Jvkn7q4NtjNx9CHZXCtYakHFE+WcOgz2FV01/IS0aBf2DBGbWsNoc9vSfrrcZ5mqX
5r1C/nu5PHXvqhP+Itdakecco9yr6wYyDlkcgOx8nsFCtTKPenuf9GSBYfrDGs+zDuoUcv82lwF8
AfuC9HUszfzfm5ZJcSGaefNXeD44gUm7aQYKBgltuybHeQUxzyqlM9NoIkpooMPkpXMT3lx9tVIb
YnjuOgMABzFHWPNz4E4jOjIZOXQQkfE+Ty+ZiZVDVcy3lbpYU38VTRT/BK9e4O2Bi8PaKx3BXgpg
mxFC2l7+Xl81eY4mAKPyzPIbySYp+6OUItkWp6aTW9TbRNrQ1vA8IV6m/vBOMJfqXd3ZIV2k+VyV
GXiJZbFKedPo8GLbf1VyqoGpSHkpCqB0yLaYCbgjknjNOz7u614RUDGrL4EcKfpxUiex7Z7gl1VH
jcgbI9wQJgAAOV6uRjy0d7CNncPnRnP0X9VtzNppV+pwWYg4O1RJeWZN1fbwnBXAMlm7/U3MGeCh
jCyfJCc6yPUKf84bD4jgpCwklT7stLI1gemOcGXVA4OI0O15levf/h5482jC8i1iRNS378fTsMD3
2vcwj1KqV5vmNKvM1loNXs/mYqoYIwPcZBLAZMjfWYkFDJoydvT8LR8UemOPzJ/B5CDCuzaNISZR
u0jGoJB/vlApMPejIGwLr3z/UqmimE92TW1orPJwI/z+r+12TdETXWf08KPOL7+ifGOzo5iR/wm4
Gcm1nulaOY0kZoC0+thoPoAM8UWScl7LpXhGKpr1PT0zbsfk5MWVR4Y85CTASgRhesptvp6CsVBZ
EKTYJW+UDSC6THvUgQEYFtwBbsTplWvWTMphOUW+r5eS/lJZRdy+bPMHF3WN3Wj2pakJtkagXp6+
g+sYQ3sza9qZzCdSmlQn8yKifkHiv9hnp7GxV+0L/7h1NiTcB/b9bsFQdX0IIQUe9smxzWMxuGPA
NPoXSeZj3EJID+kPQU2UUPHjoQfe5AuMMepraWesokqiQZfQ5p83eswsdMWcrSLvcI023vJg+/Y7
B0ouTYk4BEiDuIF3yZJkz55Zm12DrGRQujNqDIO83B1iEB1VfR6MbbUbvJcuDEemNA6qqQjOP2Zh
IONakV33s6igZjGzWLG/dVNPrzgLuKZS+QQu+S2/VQ2wbV0180G4nxAbm18AsajiygfplUPSq1Zr
0zz6PLQCYIz5QIkaO4XqOYhtsGV6CDPCSoPgvERMLUsB6mBOHeHvce6esuTlQ8mjHaTM/yJnROFq
n6jftm6IrAPz5luzofR6uUIQbHk6tK8v5h78YiRZjzO0JE5pkoZ4YQsETQatHMeXacDNk4Bvns90
w4dp2qv1O57teRRHmWHb5JkiAxLRCzn+AGXDeQOqAz80F73v9HYcH79rcIBVCFFB45LWFnSnmpXS
MctEuSRZqDvb0FXTCqQy35Na68l4XAAFZi8B+bxOr+UgbksbtCPrI8XoDi5wXIgxHs4ub3cc4e55
OQuweqY2+Q5uS8Ov/yXkxXWseRg3ja/xD4xFUjiizF3dv6HUL0BygVhWrw7KTOjz/w9ufXFHr4/5
Y6HFGbbr1KHuc6PKNet98ckK9ZJWcPuidM971g4mV1dZ2P4Pz3ZOUE9wSFkTpw0g3mCoCIvEJjXq
ZteoGazOZ6bolLC8wU/VfYddXafD4fkREZiUFnlu8HBrEGccIiEOD08rlRE9hKzttzBRowCxuSuk
7P5N3J4FYoVp+/Q13rkqSf2boIN9rNn1gSde+D4GRQtPT1ymF+4Rgp/rx86qTvuaF4EM3DGHFf/n
RCY0OwwA/+Noba0NT0ckrbr1de1egtQwf57EtH8k5WTKRrjX9w408o5PHxvuI89yoEMcOgUBcXi2
0dRoqkocZaljTy7MZA94dUcQMrqDfrCV61NxNe2S1GuQTq/VsXTqzXp2/1S6dP+m0ZyeJu8m0/TN
hO/pjkaJ03OKYEeFtljTwE5rv6PVCKGBxM9FSL08tQh/4ItQzk7s5yKgmZeBRTx0UAyLkh/Geb6W
+Qjqd1eGWcqYFR2JnFdlZOlCuCpP4EZH945m2z5YGizOlQIM6aRCRvC1JKru7OQVXXN1m08JnXPP
YSe8/f+NYGnQI1MgCBR33DJbcrXDfB550sruSE5ehdebth1sX7KR4Axlg0TtH/aO9lXzkuP/ucPv
ppIyYL7ZZiNewDVANh0LzCBDrrFiWcBqc9AcDBbzt5t7vakiJ8AS3QLY2C/KipUXzqppPqJ+XBKG
Su0iDIMfBVOe/UBVINdTxblpfpPcoZjm0kc71PZi8TI75gj5TsseRImXZ38lc+ZlgcONDM6x7KkN
ERlgdNpH/sHq1ZpeGjhAJKAkvm2z+GTQm2tVxTSDnuoPIg3kz8wSu9xYa7hTXWGG3SidJTomsoQL
Kgu3keudfjL3E5aX8y/zyWkK6CEOcwhv/+F1w4XcG95oBO9TeXeXu26j1kcrzTUTCijMGy30LwEO
yvnk+Ho2WZ24+V2ggy7qoHIHrn/9022Np8Gl+ymjw0PwDAJclpZodCMHF+zQGTA2vA3kL8cf6FIG
660aGCbVrmQdJ8ULEiaUSZ8CI2XaY6DiDScqQv1r71uwdlTf7WZE0hyv55Pe1sbv61oAkod6Ih2t
6GQ0f/KlT7GnT+gf2iYTE/Uz0+gsjvxhru/bjyqRvhJRXHanA8CXKtWqJ2ltmKUyfFTZ/hgf+duS
vhQ4qaFgiPRibHApVJHXpcd1M5atiAKD8dvamjbh/G0SQ59bLZblStkGkgcoD3/p33v7F0375pJ8
gGowXyNuWen0dNBuY6O8zsmjhy18X0yOIZUcY+1ddc2qISPx42ux1f8gPwxcQNvSMVPE0l00L3M3
+lIBNbT2m306NyqKR0HhwdLQ4+BZmPRBf+aUVcLFPYVMHaOtxixOa4OokTjGteNurk9+BaIjU8j/
X9cG9/ULBkyjkDtMcvblWe/5QsG3Ql3wjnrLTOCiTUQvoIzDRBlCOZKk47fv/hOaHNcVVkZ4ctWb
kdO+Za+O17KFeSJm17riOtpgtNKd9io0rzJmqomk6J8cOn8W6ueyT39nsJ4k2PHw3eErDUiNMPOH
4VyPps/pblA8o78NVfZTac0dDl0eD6vZ5jar8y5x0ssFbKngffhUbPfEr5mkXmU0T/zOj00Zdyf4
3eX4F2ztTn4qHR70p4z2iUzNOxhbozp2s4MpTVUDHWMjmvX1Gu3hQmJGOimSzhbERgdS/93D5Yt5
41KloM+K+nKrRK4Q9ML4nYRvU9PB5YqtbMkHleM9UYXqYyMqEucA7FPcy8MLHTIq81vt3p9d42rt
QYiwZe7WTzMLrTq5jtljE9PrSaXS15bYG8RQTMNhU3SJBIrs91/0/E8yI4A/TsgmMRzDQcI2Rq7N
u81r5+UXlk6AB+CiW65o8MqJuIntC6rt8vPRmSqb4J+k/IIAm9BtwHLq4gdRVwyw2EMs/zD2PvqI
UIH/eqnQVQfWs87VcHn5JVQ25naqUr2lr9Qk9TRi10dKY8wvtdUNaZPM0B6YB7liQ2DR7LRVs2H8
t9Jni4C3V6att817eOSthn5Bqs72mDI2mJcS248mAtHL5EuD9KXKemJa7++fIpCsVifcvq499nz2
QovHtDlqY0XtRqak/sVFGHzI2MencV1lgbzvUSrHo71d186Jm/KtSQRu2Sj2dtEKVxS3H2/+ULsY
PpP8r/5RThAXc8m1D3a7GoTSNFIG4WBENxWBu80yPI9Zz/0fgWxrP1RxFT2646INjbgsGU18jNit
VYKxn0QEEUcIczQLrqHPp7zNJuxR12qTHIizrwSS72OZ8wnwQQBnlbICgB2cN8yt76kyoC9uD4rB
+QcfOLnXFBSZ2BZDRhsDz088ttZoqd++4kp0rINZ+vpbeydDpN2lbfzasu2JTDkS/oRnd5tRPnY2
O+4S3/bHmjILlBFo0hGC0OD9UAbJyhwTcI6EYifB2XNRJ1Fdzi6k6g6ZkWpS5JxgVkU0OL24sj/a
X5RoOUccitQoVPCc8dotCaqpU95YPh2u1tp2xts+mP32ILkE5F5n9OWYMyU9Eo3YME8UhWKFjzwj
Bm3pu1S7CH4IEfnad87Msq7jq8rmC75ofKqfhHRoTDrLCc0f1qu8AQBrgi24/u/BrSFTwch4cT9p
PXkxiguFLCkCE6VHkh2SqKMOw3AsjPUKFbO01sND/uBXmWyVjEb+NT+qWQ8qcQAMvIEsEJANFcmo
C3IIQsrlYqqH+nlDjMX9hUUkNI51dHhtKMZbLTC5/5QZLwwNNTcPWWdPLQhohTWlRm2j1gQ3DrVl
7/p/YNscMkAC5GdOsDo+8FVWIeJF1yz/SwKs2JEi3ksE/v45ygOihrrkVX8TtX2D/qf16/LvetNh
Wr0o764q7CcGc381wGmz3gwS5Et5NnIXTnE3j2wRtuhlYboJoh1q/fkb0tTXHaLlsTgJ+2sxfIxq
0d+2N9dGXuZ4bd7+VEUxEmz99/uUpYfK65iJuFfSivOJ8JNi3A7I7DkA6v53ii5eWppz1i9UMe5E
veCtUnMoht9VnJFQ8NK/nAkhNKBqnvoqNouAe/LpS0ogWDHORSkftTgB71Gjw4OLYISa17K4Az4p
uWWO63ftkQp3d6AOJ2i5tqIN32Wjap7PlDbDcZTs8muhwgewaRki7gWXNvtUYOrOdn5qUNOElo1B
ZfRHuX2DqbDQreSU2VqveV+nx8dnmTmau3FSfV7oMdKlMWmpD++yUASQo4Zmkosh+d1izKOQ8VKg
6puTOMS/HZGEFwZCPYFMWyzwB4j1+k4yTuGnZceq5AAzUhBeOlYMTTrtZsi64IvFOWMScm3T7O90
4HRqtO+hHhoXgr3ssIN32PEPovl5YeWMGtzmm/p124lCSCloalLPegIEDKZ+pbhn0kiKiafWBYah
+rjcvo7F/xQC+R2YCO8/A4CqIvO9/T5KJ7CgZSaBXtj1+m+jzjg+nKg4kpP53I32c4NwKiq+DvId
/ecWBiHvIuVlMyMPYsxEO4qIqmTqe0Ox8IVcyX/Xu/0YOaCSXoEricnvPQNNNy2OOpP9dKRlGag0
7OWwB9BQibecr+GQ53VbpbtBSYW92JjujluRtnegXANQQiwGGEFlSvLWvOXau/XSMq23hU4ywoTw
wEVo3WM/gOJt7kSfr443jS9RJV4Hehg4o024XKtDdxo8kLOtOGHovrHbJv/IgT2RWxowvHNYaHtG
UBI6WzuTWYJPJx3uOHqRtDlsxD4W+V9kiCn+3+U1iUwdFa545E+M456LwaTeS+Gv+7NiXSqgXqDu
X+t0zvkqHNkkudiLSSItYT4cQJkT7iPlLcBOi03bUoivLYsMYyneL5YgVlocJ9uoekra6tg1i1HA
bT0e54uyR3bcU89wEFH1P71SQR4kCfEn/gtGukoqb1qm3sZdy0lTK0jxUOO+mxu52H8zokdp2Xal
/Giw96M641g92aBBnK/ncbW2Zw3CCBP9QrLfP9BdjDDK3RsMwf5OK5mq6RB+zbDyFNl+0mNU4FI1
+p5i7pidK5WlYcawoJn9lnkoUztK2z9BflwfYqtqXRli87vPpvS1LYJP5F1JJ1eWB+H2/8mL0tAr
XH0+vuWmqNpu8GDUIjc1M9COVv6oz1Hy5bpVKlwXT8l6obfM/Vqe5O4t9q6smM2WxedN9UU7KNEU
3zKJ7HJaB5/LfDlSWB8ErMs+NhKrT0sJNhqWNiWnkHLpAHaNV/Ss3kcVSNU3sHQpdYp11c/GCvFH
IxGc6dnIjgndAM836x2NLsVjHBt+gTv8aC2E3mbMBs26PYiSOrxtBGleJ0f/yoI9MF4JrkMPY3Iz
6dV/UUT6W6maQorFd8QDqTHHT4AVPoGgeP/TUQ6nkV/DqGxUtJCrf6Ec47LEUxabOEWL9ZLzJLiu
IBDDg9JcPsUCNu12ergKGXKkvX2fnk+/obDdHZTmvuTtKTYz+r3W1UFL92LZuuUZC2jUcznY03dk
ubyfkgK1DdWziLD69sqy2WTuZOQ9GZB0n9ALAbu4uBO47nvcMpAOPSBsg37raE+0SxVSTaLcPTtM
aXc9BCeLoYFu2UScB7t7RF9AR4rgO19e6s4uWhbck5SGgjicWKjChxwNnog9+m4MsbeVSt3rFKhA
42fNBCkePCSU8iEHohiH09bKyi+5qMKHK80F+DX7HTI2DlmAvemoHVxN9P57aNrprS3IBtyzN4uB
jbeClMrGHg3LPQoC6xtOIgvsm0nkgPj7U8c6uUBb+DVFaC2Fdg66AAh7c1APXEaeFm7FdD39NRWg
IkguYtg9OijfhzcemSTEwHsnaj1mZiI4TtELPMGAuHMS4UGSeyaVL1RnOVUKHmFPurbBljk9EU8T
ncoAJi8OZpu1cHZPkEjwU43EELdgX+DTnLGD4Na85uNEUrKvRK6Nce1Pa4pyYsgPk/oxshJ4RoVA
nbf17t9x4SFnZ1+D1bc44CllgASd8dsdaHLyZEYkgIFULP4e5fE3gGEOaxaAn0Y2F4TtHhPi8Fka
E9HmJW1mB4SVKc7c3BLj/5RZT5xL+hlM+Z34uCREEzR2ufn9FXariauYI+743JRMjPxvx2zqOKn4
XDtdtITZ2ITksOt9AvZLcEwxzsErgnY+HW3rUit9UzKQIrVgYTePETrEV+8eRyF2Q2F4Pq+qZZAa
L5dWsSFn+t6D6Tq0BDurvepwu7Sx3WxHn05NDwmwvviF1bmdH6T/K8GqKoNdRmpmYAtAvAKyITwO
upLrrlABfcOqhDBZYdgQIEIT6sOQ7lUrNd54WF8OEPlFkChXhAGnbNEAkeUc46kol42X42lOF0Ea
iwXiNLbJ6qz3Eaehz8Gc34ryqZcdPYbzYsG0/PkAM8eNlZJPfO35NQk62nuyKBejHUakjYhikeOq
cicByc5ZbeLOfkk6Mvl9JJbryJf0He8ErTY7nnoSrvktCPGXpf0pxHPxWLe57Ywfo+tqRwfBKLgP
f9fa2Hr9JuU4dwt2Xa3zej9EeWX3NkeezrSA+yVP/DjDH3yqpEkx1UBDFC2xcqYd3MRV40aJGGeQ
O6Bu5p1t/XcKOxMl7MoEvz1jQFQOEr/gmDZ6wgeLEW51wE1CTuxUzetGxJBEb7LWuQ2LJhy0V8iz
s4QBk55lKFiYSv+Yz9qkxGSBqd2naPBWjJU/FhJA1wAUzQKV2ObOiu5DzThCbF6riL6Ej9sAWbSR
O3oCjBa1f1f8TXMdbGv3oKl01AsZYIf2vysweA9Ce2pYtgVR5465eR2i/r1TNcD8ZUxD3Xy12U+F
gxKTTWDB0Ck6n+uJGV6DWWHtSs9AmnnFKxe2PpZMbzQhhSJKCd7SnhO4vCqWfu34iXTQ5kHmb4TL
YwxhCISdKL+K0WWIXsWZ/SYebXGad4tVhRZ5nKFBlW8ORf878oNPS98jkjrIqJF/dGYGnFXMCyRN
wBcjn3XbsgNdGP3VA5aDPp/xdjSUZUqwwuOiezdsFmV2xrl2VUei52XRpiKnUhjF5WpwF9K2oCov
gUFPzCuubjBEI68IP73/h9clMWLAzMUPDYMLkgeNeYA1cskK84kxz5wfhA/JzbkAsOeQpmumamAt
fc7Nt5r4JXT5ph02y8orsV6kY2Ha0dioLWZITLvaSQKu5vqa4X2qv9X/IsiUyT2KtBBwNY9IS8gv
J5KDI6+tETVbWYHaTSWAkkk8spZ86RHS79CB0sxdmsjNdRbZJV8DuZTYJScBmnbYIsXvTkni6+Yd
Hs3woH/9SaUmb0VDoasPPLcn+XhDDoaCcRRKa/N9cO7uDtk9GPvfNFpH+uk5XrtbJQSSQWwwxLos
IycrUMUPR9CECZscOHttYFogO4SL9fGOskXhjvwGg6OxwxbJf//FMJAmsD6xc9WJFJ3wXe1UNBfM
9LEIDuFvAymAfvu5mb+9iJk1R+Zx8gjnlGIogoA6553iY7Dft7GVemxm3NZvwy0e6dRB2TwRbPIA
Bi64AytqbQwKh6S4cxvdDLYC/6+0212VOiI3XIpipNcZ/mopq4ZZ4CWK0EENjaKqPTEuB6slTpnP
Wgcd+2YkMWuUcONvUp+Dz4BovpLHSgZKP2X+CM9mqj4QI4Fwb08EiqJSkx2W1uXXlcO52L0i+ntr
9Q2Q5DwJThuX/3uhpaATRCJS11e+OnPnKTrgjDjGuHQEssCAbv9B1OXm03ONBUlE7M5DkmokZafy
ipkhDmG0sTnbCK2Gs8DFYr+Y5El7hUEJQx72ff4afX16mEAaGLlAOFIDniC0l/p1ZsOcVRpi4vtL
VCO8TbJXS2oFY6jkIzpSEOatXai/xzmbSUcjlevVXfwoTv6JZKVW5KzFcSXkzrJnRRILWLihvUWv
1AF99k5Shr7SsA7bAvtYhXB31wjn9sf8u7tvLWBrgChaiImrBVKFydv6DLFxjB/F/b4v/BsDhjDA
tQnqu0u46emGdxxZzGK2xfZfUhTRkc02QYfWjGZXIUfa+yjeR1QBZLRIWjKxH++5f7DLhxWiFzRD
An9glPae6KAAQC1SkvQXtdC6O5W96BTe54/7VchEdCnNR/aNJSAz+fp922klAqdDVoE8b7m2taFL
8Y7epG6muh9nO6Eq0nEGPE3njIKjlRUkON1Q+euziLD0rGNAEoYIKlvW82wnEFxWsnyzWSCmfkpJ
3Ne/nchjiPNffww5A2kgfrz1db2UNZl1TX3GPhFH9+p/O/vPBCuFcaWeldMS1hgmnGsPdGrdKDEB
OF8/RU3CSTthwhEi/X55/c6sEzI9mFoFCh3LXUSNNHfxx3CmhPVgujgwo/p85YnmHRjkxGPl4WTC
x+w9XqmuQXJDIrZfKTmxim59m/A81lItdmlmTBsOPSaqQpGPac23uIL2uMFWg5nAgDMJx8eTjUwG
OtD/HySD+9htUquy3wkXUp+YfsweVGXviXUiuAOLBDipOWoJlRXlF/Pqozhc1Kvew5YcgnGb8dWh
mFEk3Yh1MPBjfDu69XvTyhK94NPhOFZ2pZ5c9xJpd+MlLppOaK5BaIzlNSBpduJU7HddM4eaLzYs
PkbX6z/ljYK3gF4EWXoAIY7e8qbqgFylr4titg68EBm+DKQD3my0wBvzOuGJIK2o3khqfbzIyYLN
NtDX+qO2ELo2cIB0g4FmZtpiVfeD+3N6ulYhQicYn5GKP9nR3BW9vXjQSAAnJ/EYGFDw/nVtR52o
qeWxTCaeRYGvfZZejeEf27xOYMW9dOhRlIjd+6dTOpK+r6e4aYkKarfv37uvswK9ieELzCJvy6VH
u92IZAjx6jsqFgFdwFJn0KDFpD9sNvsnfqyeSFAxQjzeaaguDDzIInvgNZ8NHL69b1IaAmOVFlJQ
wex23QqC5GfEmBpZJ8//fQQEhw3WOSNkJzFawJFRa+vG4X4RpDNxdnrqLgUi6t1H0cawbYwK9Goi
Ic5tL1kxi/RP8eMp6wsY9x9IO7PQx/D0fyvuVm6ktzkuAi0djc/HLq52/E+fm+jz5foaClFH/+XL
31OsKB2IRsnvGMfe2ZyxgYjZPTUeGnObEOcGXI2sHQIoG5DdopJRlb/rLM3rLPiNwvBs6/4AqGMs
aQ2JIH5Kp+VPanLZsk4PIlEOIpu5f9BwvAZysob2t25CktSAQkvQQrNfEVaZw79jyq9nfYDRfD4Y
31wP/wj2dpj8sA/Q0hr/mxqIp2mF1Xvl1WAVKbk5VGmJFr+hGdM3Ueq+Pmcg63cSLEnCoY86vtRf
4Lmx+nx5Y/INTLgvJKteSZ0Eg3rSFNWYVphZEftABICjkthomnBA0L8AkM/dzwRXKWhGVl1LWws/
SY61TAE0mFETK/ISE+xHEXx1yVtcQIpvtTYYez+Rw44aWMT/l0fPllGGjajOO+17ExsU7VBGcDgA
3yldSYsMrMNwZxhMOQlGcdzlcjBkTqi/yosegKsKQ05dHy12lHUsCq/oS3vjQkzTz2Q5DcJU6me+
R1wGoRm2xvevZPjPc4Qk+iHD3KxLGM6/fgtgRPJMD3/dLcRiAOt/u8ROtO5I+LkOZksxHPTWksmb
hYdjH/7bCUAg18bNKN36CAeFzoigp7KPoL2ykiGa454LExEq4CkZVyUNuxb+AA5KbQ/hSL64F5K3
kVLFquj+qhk20d4NxJYxeazw9cleE8BGmkm7IOm9tPAQDmCX5shT0n2fUPsWy2UqBldsv65szHOy
vsLXJkigF/wsIe5jaieghp/xYdECj+I/sFm5x1QkxopCD90jLpHpF91CQ8GmRrRhQaAWRmU4BI7x
Mxzql0sgsWWLh77xihgEV5YxEV1HektB3VuyKVXNjAN7i9iOI2ye+ogoJ1jYOGirRnLXtb71Bxyy
ZQd3dAYcNZRS93YnuvpxXPYw8FbFE1CbdTXDF4zbNLWavJ1AlUANX710LxjkiQOfJ2bYdMq1ePuc
B9TQtIsUIWOcMF5gJMnW5RM0xCu40BWFH/7qjq1y04n8Y3FIniGcrQ4Vp7WwMRqHJ/4eDJfmjSL9
TMaFIcqMTZzHXc3h+WF/opRmoJjxU9Gr2fJ5uWRlBtFeAzxVBkE5onKXrmLRmqXdPIKVBS0GDmky
5bd2m/Mj4nnCEIIZ3iSNm50sU6smJuvA/ecY/ytZM34ZmyicSBY0nm0qRbDAAjzpmDXLN51NowVY
+MRyHP+QmtKO1Ig0u1lYk2bK+ZrIK9Wlcd/JpJ3nFhM5ykSllzKdJiWFTvEisQYpww3epvBEqqRA
tFBKwXxIf4ZMFunnJCpRuCJUXGRyx/leTXfm77+rIQKPMb9I/q8U8Cy3jIik/vEEzAK9VHg9RhBb
0lxjqYnhfefk0w02KZwpOP89jKKdgMYYt/xXPtyVmWDXCNED4UyFva7uDU/RZ4WtZ8aXw2M4AvxN
qb/ewwYvtl2DQ1YZ/VT+l9jn1uw0zLDMcDh/xj02v4FQouk7waeI7rSe+aNOnn1QCaAR89EG9DVl
zSPb31CAuQSgajLO+UutqP48wz+hK6y0xqY9uVGiMJYcbsWevInFCJOMOYdwZ3E72rSupDWSORSw
zKt/haKTgagYY+6wPzIXDNAoPkqU0aPioSlXv4GM6WGBMa4XbdH+Rf0YUS8Nc+vvBewKjSyRl90x
DmT8iB9Tb+/KdhWOAjxVcnqlu0KB+xjMLmyBwj/qHkq1zInLhgLHeUWKBONSeitThB81fVGI5ZIK
5dMYG/CYUSVlhErZhAzZ9j+qgXU9WC8ReTYroGXl/UNjxoRdqQ4ohLTal6HCf+VKuu+uzrCk9tl3
SV5LZoivoyS6x+gwmsEKPkUlVE2abLqqA0soq/S7+/noqz1jNldhfeI3KySnBVAuvwDXICAn9yBz
JrV7s5QpNmWAUUhXGhQoy7IoKkrSP7QZEgzl09phFd3oglU8IkJxPAFujkKvH1HLNdmMnHxYGuOf
9MIzT7PT6S/m4QsSiBBX1albprGRBuS8SnVy+5kliEDktpGO8ut5R4Oe+5BAVPzyP0AIw/2BghEj
+86Fw49EPpGCe7jvrtlJtJ7ZVXYziUBhMVoBVhvt5iIRCq7gui5HyzTVg8yS+cbmK7Fyyn+EH9D8
KTiLOoZilHdP/U+gpX8SHENPoAdLNfFum9m/dIbOQ6ZpRuM8kP8aOgOBDVQOMygpUkMRGXdOI+Fz
951aBvATy9pYy/mp6Gu0FNa/ehbGkTLUrQAOL1o5uVqTB0K+Bg+bVIA7kZOOhhTYToIpKus8LZSm
CpBcN4D6hsKIgw28se5+Ae+kd9lJhNsUitROooZBtxv4BHcgzGN47FYvp+zpucMrGCOKZP2jnNpJ
rKlXHO/Y2dhiK2g7w/ApXm7kMvnG/2nkdn44BMk4/ZDLbd/ECtPS409LKqXpLP1tXD8yUqS2bwtg
m3aCHBKHoxKBcRwBZTciAlkd0tUhQ+ryEQvPzUKWZeWGZqcv2z8MFY5fnOJNXfjdtPHuDhPADBop
Z/IvkaTRUsbO+Y6GmMO2vDw/gE1YJdgxg3d7VWWneJXMCMI5K3472YhXJhW6GnplXA+npkDwREqE
xNkD1mrJAXWenmxDyhlXRNp2xonAhLg30v1llzAsZ0raXmFGbYFDmT0K1Y6yvFGt9m425W2JJlON
1TwtpM8cY2HWM1y5LO9jfGgzAE1RNSjaOuK4FxqoBQdCZ4sAS0AiFvJGJl/55FUwJlmkzxqUzVvp
N/2yRScOGJx4CbUxnLmRaRb7kE0hs+G+I07z/96nhrRRegOOVRgqt9aiD/LmBqNl+YZpg/YDyvRS
xwQh7nZ3CR2kFV+qO6AEzwTinpGI04cvy8UpRPrQ1GQKTt1sp7ZcOCWwWTFyTKsm5fjY6ikyz4aL
HGN0VuSTHUwtPQ/5hzLayPAnwbzyVepC6JjrQuQ9cJUCtijEv/5wGAorcO9ZPBRf+FpMd2LAbujI
gE6TxH5x2qp/A4HTiOxnVk65znW9+fWyNGbda5hjnS6LejHwTlt7fBz9smxGCG1fa4n0jOWhEUXn
kDoVW7e3HbWPAVWKPL9ZJi2zpaxz2s6+ZvfZ3WVemHMZR/7dESovqiVE0BpBMG7IhBItvuxkhC1e
18y0y/pVA/EMTSW/Q5R3p+xi0HHAc6U7kwolO90EsvRJctVLOJO2VMGnSmQypxvFF0emuldasY1m
0H9ClNewseM1M787D1OdHGBY+WUiPl29DL4IEbQ32GgaRkcnWBijb51mJAbUqtGhmRxieyCF9Dha
hqCKoRjH2bTkogp1UDELr/e/h4bKzXRTJecHdx/GSLLkjxVr/XwzA/3B1u24WCGfBLwXI9/RKeQn
Vcq5CUSJQMqWKB2XUsCJumiKxYPOGiMKbFYdPxnsNecJmJSy17a1z1Z+XljoORPzggH4LdpTzamf
KiKy16TTH0khegLmdv1hfbsza3BOTUmNB8ZxaSCGJQYkiI584xu8vvm2S882EhkUuBkkN3ncNld1
qgy/n2kYaAS7W67eh+SU1xpK3TDK19LdUwFSQo4BZ4YooS/rF+uURncgIhujxFb0BtGz5vUuIPSL
sdQj9ssIWRCe/MO7f94B/REux+hzJmeSCcDqKzk4OuxP+NtGLWPbybHNXshEbK3CYQOAz6Qoyfsy
YC+7yYM0VR63wszacDDoL4ekQL7RhaV2m5MUWWAUSYdIl4LcbD0S1n60iYBQCXRyyJdF1tMMuypG
1UPQSK3W7jVtU7JcOjKUJuL0a6ZzJKapNQ1ontR0HYPvCEkI5Cky4qRb7gBj82NdtCfOKmfRu2nM
w3yOhURmLCkaZxv8zRuhvPO6xUrCDeipYTU/RRpc+O2O2tc1RGAyRFNGtqPW4yf/pmqGzFUGRhfY
4XrJnunhBLWyTNdest9UaKTr9dP130A4/ENcVIB6AjMzX/wMxDmCwridqojrgIiWRdHdzuDo6KDp
INzLdWtDRa3rcecnCGUAucPEJdHKC6AD7U0h7nYApJ71nvq27AwWYQqnLevU1I/QH4yyIhq0W65/
xzs+FWJCRIjQcOfmslJbunVgrghhIk9DC5Pr9Fnicx21U8myWr86v/TdSXm8yFx9M6tIwt70aBX3
OvCt572ALf/YKF8cXlE1nd4DqDuZczT4Ksqkxg2n2LzAoS/zanAVVXRDj4H+xMsiVV4r4vapx0L8
3+4tytS0wMYrfm3T4t93SzT0mO5cmsMgcIGg6jXiCb+/TyvZDUuFbfqSEinK/UTH0HKRD6HpqGaQ
OgJuql5cMawW73dvABaAM62UlzA7rs7QaLew1aaOq46mBNmtKiZZxTSVU1GFfH8cWiqqvCHGtAHJ
hJOxVzGxXecIxqvILPRpc3M1KwmS25yu+TGF6BHfSilbagmhJahgzqI1HxRD6PuZul8dpa4ITrmZ
opDsCgTjC+gpnChaUCAPjFeyB8JUAR0uk5IpNIJSJtSpdj5fTzVLPETMhei9t5aQ1O5RQQMsCZy1
nh447HZTYtr1W7QI0aSmtD7rRyr6QeeyUqtdKWM0oWhLRB61DDiC85aXCp4excwM9vrFGSH+BKYI
Gqd7pRM4bqXQ6a2PXYRsK26Rw4oZsPgwEiE0t2fjlL8PapL4TZ6EXQBq3y7+GzBujVUMGP1Epx//
g0+3uiEdlFYhP+A8tu2PGl6BgrSIZZD3JZb/rupOLeqYI9DvSFeMi/3aXSD5etowE8ibTF39F92w
TZksovGo3jBeXPcFmBhtGhM7Bck4vWnVCs786PbaRepsRAGyCfVGncVzSBK3pzwuODi9MzPyxrkR
UwqL7bEFpxfUlWOb+7z051FiT2SMYHsq229hdSp7paXFqLAtZs6e8hF7AukZDP/0LDCObNjWsYTN
CVb+j2LWQLdZ8KayxtkcvnLlUbKEJ4Zx41LoJgzoK17R2NyhgwF1I/jcvCGESnbtCT5Ar2b1z1kB
tGpYa91aeIzNP/pCVekMhC3UnoNng1sNSOJh6kWHq05RpLmLuSeKjy8yjxjKF6ud3hOCFteFFAUK
wbiAMO5CvtJoLeOvIdniXwdx6FHcVTcfYsH2aZfi2opfveXaDAYRbgNYHPxEvBI2XBHGD/V5bSAF
8oBA3vD0KXryQ/EHx5B7SGyX/UhinL2UAgCSwQHVI7H2D013hrQngj9SeWF6gJNyhF8UmBQ7kFv9
obRb5Ll05q6D88g9WXXqtkbGSrgxKBbN8PpQiugZddGA63s8TunE1P08cAAS40tSdW6/IjPr8RwC
oNWwU1rf7qBP5pca83tikmK3IMmG9xKRLepW1q4pnwkADEu3Lijv6yrVwDJYJDYvfslao7FffnQ1
K3os6qFIxmx09GayXAo1H9oEhAMS1tcJ67VCGfMLtEaCM/wgtAafd03E/daVbYGVuUpCTl8FeniS
iR5pw2elG7LY5XQdwSwAx5EDWej9WHeVuMVZJ3oF5toGQN25HvuHmgf1YZsfvYdAktF1ySuHJ9mY
o6lwnPovvNFA4iL6wUekV+k94gL59+Sv/EoeRWrI1t1cj5gP5kJ2PpOTscqkvHN8tFR2Pb4mp3eI
zl1A7HG6XXtnORsMOrErsUbLQtmRFmkGs0XvcMihECkXoNGNLqq7O596/7fNrRQfvQFlUgn6/vzJ
R1ygbeTcU4JT7wrbgJLX725gIPYoIsNHOoRlPv5Wv8n02sIvw9MTl/eRh8/mvORzAKnC+C1zhK7W
Zul9nCa815M/65yAI62T6BuhrKhWntYNTNakQV0rkEs6iHBkv/D7yI3+llvFF6BynXkwsl80PMDV
tKnydHlFInphpvfx7/KQ5Dn4qPeuKi3DiVmr6AMHOSo1N878wJLCo7bZWVVN3/sUWZ2/D9a32VJA
MC9lgy/FfAf9LnVRxQDIB/1xRXQCnd3+OrMLimSlGKl2UJY4sfhUbtki635mNILkIsJfZMn3EApv
KcexPLzn7yjnBhsK2FP4WBUwBTj6UzNaNKIugID5Fqf6DtJu+CAWiTo5Vs8RrFYGcmwo79wIntfN
doTFlQpammFd1mfHIDhZPC68wEsHyZK4+tYbQz7pufxNJNgvY+781bsrjPSeylsihnEAN3+mAb+N
NlKn8MUE1bHl/FlpVdb5iQqp50cYQcsPdDVYja1HtoOVmm69jtJ3hrlgfUy7NvcGtF62Ln1/hnOz
yQKHDTb0lgVJQnI9nhuJdW1SOR8Yq20TRWZ9s08pNH/2gojnXNOntBYKSGRsUtJaTZuSlsCdqnDK
YRz50VldwiQbASzIWCzoOroNbxswBw0i40W+wpqvNpUl3VjfYKSWxJpSZHcxI+EspTuavbq9/FWA
iV6XLmAv60kM1tis0vBtVg2TRJLXeS7zRPwBxkI77nGikbydrN+Pi0e1WF+sc/o/4ugsI8FXoW4M
eJsuG08UxppP2hDXjDTMKiANaq1wDwPnAscfUC7QeFaRqF5/QiIhwlW+vkeyHCE7vCQRPkx9PZH5
neWhupdETimjMD/wSiPl+v2PTCz3yHi9X/w832Uj97pgC+CfktjqluB4cHw39SrCnqrE4ytaAVcR
Gf6BuOI9/gh1ZaQ2V5iG6sR4XvK7sF5/GS/xPS9DniXiLwFYKnRSfR9tNGmYaKSf0lvMPeT2vj0m
5szouLkw6l1p/1NA8SuFj8pPMSWq4J/sBC8hkHw8GT5tO8TawwroUzN1scCt5NzeVBGosfe3Ju1a
7f8AD1ELwxCdW4caePSRgRpPUhUehxBY5EhFkbefhi2zp+9F+PY5XDth4nIee0GxFJAS564yq2rO
D6vok2d3WhA30fjAxEyeeueI9V2tHO/9TUdZ5R+5zXjnj4clRAOBXofLQAXaFl0TztmSDLnpr9yP
JHWfBN/VuQ5J7MZMLJ69LrI5UZfwHZq666Hcb+wM4Rz3carhlSGKWJxq89meJeAoO2kuX1HAuY6a
OG2MrtUMTk98kCoNgQUlUUvg2CFXP2R3TlgXMw48V++4n5cauWq6PRQ+8OhSsh1DxH40lLrrFFa1
bc+Ipa8b8RVQJtnmQLdrVxoxt5imdB48Mi+jI+aJa/HCS/Wz1seT0cX+IsAIxTXFnpVmIrTeQjX1
IcwYwf+Va9sdCQdVVhrFsl0kg00trtP38ictV1qID3t4FO/KUu0dTOnGaK8ap9SXls4Xcq93O7E9
2X9wf8D2cat8Shw4EB2Z6A3TC7GeETuqOwvRMjpN8DDU9g1X/Vm5eK2k19+hOUNk/x4XNoRcnwxX
SYFJ55DOdlk2P+ya9EXlv1faPw6hUKl+fVBXcKuL838Z29thUXo2h+lD8ccsybjPMcxOEwtkP7LJ
82OxC/0fr9iSifqTN94fR6Ob/fCWSZZZuymD1peEZ/VF/EWONLCaGR2gZMZOQ5jEze3myuksIiXz
mKZ4QMAvKcvz/0Cgz3tG70wSlkyQZbU/yZMyfh+R/AVoALwmbJXiLlDL6BnwO+40b/VAzbx/cxhX
YmMT7KJyUqeKLvbJRcXx87geTDV7dHpwB4Fz84QOuQ9JJw1cEM2D/gsF7ez63DTFhrkrqtdP3rUF
YnaYfrXlAg0PjC0u+Yxx0K9ZvKDYwphoPSXHTPIC2YtdhdbHHQGa/QeKKd2Os0ex/TQOrMG0CpJp
LRroBlfHZzMMTNa3hTFByxCdRC77p7vbtqabQL2seh6xWLrqBUhjkC0iC+5uLCtu2zQpYK0m7ruR
t2sttWw8CmtRPwMv45J8gwN2In5wLl9FPq/sxc5UB177oOZPGao0eKQEgSWIvHexQhVyqk5wDywd
s91/Z4aFaQAMLfnisJD7pQl58U8xTKQK3nIw1F2zCrdgb/Z//gfzFIG3WBfzxgxMcb//JCI/1989
tiVM6r3IMl+tZ1aGuY1I10QMR/PyUxc64nQdOJOuhtle11+I70d8mPMLL6yD68qAUFJPweGjr3J9
4xWSyFdYSLBS97ZN313pvzY0FLkcaqiNuoI1ORtNMsonHe83U1x9Ecn/ECI/ZTHA+7RU+3Se3cZx
0AbsHq6iMuhGmur0Jd7sJAQhnragHFtihYKWWB7/C/9FIh5L1LNjQKup7ssEZ1pET1G9gZ77iwR7
sj1RKY9j9yhe6TXTvfvfgZjfJFIACqkbXQbaOegq8denU+IrdSBRbk1wx7c+IqJHdQYtZjgUXCwc
jEQ0d3tpVPhfb82hVqe4ZT19Zgw+t4GMwsGnZf+uAKqAbuwiAHGNNGdMQLV1QrmDwwi+DQf3hJJc
4Zr+iOmtzFnWonNDmpmfrCoLmqbsOIrOzRgqslWJ4kI0N9kyEgaO9FMw8EInRxd2vOE2mBawO0cO
tAm2L2Rj7YWVbwQl2ll5BEeualA0DhfXg1J0E+E8gGE1QN57di7jcAvdjpoMDtlog+Lyu9/AI/t7
pABP4JJ3IyyuK67pOy4udAxtnUGhJNIjqwKWQKAv8GupksdYFK6FTFTALDKwIUxBaRfpecrxKWK8
uHZqfAliSJHZMA16RBJl0aAyjQEHq3MN+TJ1jP5OIP9CM1Y7bYS4qaFU/baaEfWLRwBsEgehf9wy
cMNCcNAKFVAIT/PmTT73WkwpsEjptmZonpUmAtbTpdZaCTYi8A3WJuUNaUnL6mw2S0aPMM3t9q8M
MD3HpnXa2QWV+Ws3wy7FIwIZG/HFAvT2BljQ/hM73jqHOnqXfOUQi2VdU6vH9Z6deAmOko/O+W5D
OE3tef0uXvf9egfoIiLwlVTDVFwuhxqlxwD+ZAy3D59yAM1UXFQ8/a66U1qdChh1ue3Wx/XvjV1m
9Rs/hMGymy88prwH8qo0otVj2bSIQTzczA8f8UuLUEu5r8dpwUMZA9yE+2dH3s2Pf4lbKg/7t7rC
nELpjqR4LdLmVixIn1vdTyfd6o96KerZOls5H4RAgJog8e3qTFzlAj6/l6mJb+k3kSPIUxNMLZhy
4AGSv2LN9miHTu+KW2iIXeIqmrAS1jjalD0Hj2J3Bn6cjO63iwOa7Zivcz9nX2cum8O7Ok9mOYUR
MWRcM21mJcRHtkEyUMcp0q4EiEYNihWECFlwCILFqxGbR5w0v1o5Z7n1fBB86Zxh0QwD4oKA1hkw
TSeQnOx6/14Oo9l4kUV9kSKMSl68xgEpq/mgm09I9uLkn3CPAu6gOI0YcjwAoYVIymeZ3Pm/Bv+8
A6P1jpcMnzFZg6pSZFASJ6KyqaoCG/J3T6Ur5YCkhAuVE+D59cr96JPQYAe3+tfo8qtiWoh3gpQt
J2GwdT/oKCXE7fCznZJs48laOs5YwtG8/PNFO4BfFjUCY2XhpelzO7JfrRSEKD8jZTL5A6MCMfMP
iACKuxSbNWhS5ROBk9HV8U0Tt5G8nx7pm/op9ECCvtoZSGs6wFZEoWEFonXmq2+MESeeRRzEexYP
TODV0GA9wU+kf/HD6l/Hv6gc5Wk0VVM+eQJyTI53HySlvuY1FkOFuagvw0P8sH5aq0KjCSbKJm1J
72J0c8zuoIIEdnkSPsj/fUPIdVflMGIPRxQDSCr2m25gw44kD1X/S1y6OBa19ovp+4MQYuhATUfs
xzmRoWExrEM2NfVGN3VDcboMJs9G+pO1jgN12safvE6Ahw49tdNcdlxzq71jQJoaIVKXLipyw0KA
dZVUukjNFNfQfTqJjM7/J1iIPvnjVXaN1pEkYIA9K1/Bo/P4r1KcpzDOUXxZt42esI7QmYvHaRtA
qvfWA9bhrUygJw+fQ9U4CeTB9OWVeD0waKHW7H2eRGs8KTP9VkYRZJrNK0aqsd4hjx4Jr6NseK+I
i5mHN+Ql7slROmIP1gqVQLtJtDZRjOf4CSC/tBH+KiGq9KsQ4BSgN0HdM3BbhseFhPYAzg89n9Ql
jsQ2erHKLd7B2G6uL6cNAqPDkAqv4l4YnknvK8QkxOEs9iQJ77DK9ycik1J91WE1KksDYgn6OhvG
b4SuieMwhlfco615Q8yY8kvs4EFAYvln2dMmRINQv3d1HA4RKigMHCjWY/j7+OTTO2i8S1sqmjU/
ZJ4NJP1wVk9eXwKP35EpIFv+E2I4tk/BKViB6yaLruH/2E5ySFtC3V+a7SnF6VT2tw8tv74WcFhp
NssBBUYXh9Jijh2HzF0cofOFv49b3YS05Sox9OqxYUZIvW0OlwZc+p9/3beJd3YJnuSfqrzndwk9
oB/LpzvpfvjQ0FKvZD9Wo/FMDQFomfw5vrSryHfpOUhsSk/WM0ch1tNGigjEpH1UotAh0K6gosOY
uODUY825juZanGC3jbPNWOj3sUDuTRg850PtY+nfUYWVmHT/2aia70jVCdTm9qw7hVb7nTP7i04L
/tkAuS7+wsiuT50c1XgA4WNTjZRg7fXzIifvITOIQ7X+zflTeYI/ONFFN7Ros6dqQqkLOLPAMXRF
GZMBRV4ix3Kwp2E219FcxINKdF4TTVA2e6zcBZN/u5+lh+AgrEDvmmazspmQ3zEMrcA5pvGs/Xeb
PGPDVADlKb+AmEKK9/yvq1lBtnML+fwTyu9/PtnYt2GJTKvjXsUgdLD7P/t3Nog3llSEyZ7R5cne
E2cYl/gP3vtVwuIFe3du8Ae5O72W2yHDuZEoUkDsv9b1eBQ795Q7P9FUz563zXwHhFIqrnYIH0D5
lerehB4jQrbuNLore0hZJ9oyMkWRJKETsPdcDmx54r0LYR4QfsUln1gOuKOsCzLhBblJBT0vCAuG
rHEZMz03TvKyY1ePJjsMHfUxrPTSsnAd9lS7eBfsLjO8hC7yqu7KY9M1Q3IorPd09GApLuZjdrF8
4EkCV5dsv8hZsYFR+yW4kZLr3L76ZTvW9a3nxuJEZ/fufWaMs1BAUzeVnyCvZG//c3GF/bqcCDeC
XtY0Tj8gxUpNy3Tr0FpOUQgFaGTfk+ApL4aeyi+Ip0EzLs1u9LJ8tp0k+PowoDTJ2ji7+IGXkKMU
DOtFnuQHQIvnSa/OMZxQ1qwRE9usYoV6xPH68RHzklWA78GCeYlfrvUH4DdnkC9clRqSZYzKgHFo
7n5J5ZYgs1q5dvGRS/cfS5Z+hwzJI9q3XI+EijghYszvNqS+91luofMsyToA3uOSMzUHSz+uVr6k
g76egYC9pc5ORse99GNBR3XTeOuP9EJOE9dhxU0fvQMI4kxatHt37AMVAJT+J3+i9gHFJ0VZ7rnS
jwqKGG+KdeGotOgpNuxyCeunJ5pqQ2rgskGVqt7ynUGiQbbRNHZTTINRRKGbewGwEUz18JQjiNCo
v/UZOv9v2z5W2cYCEYWfSAkhZYgd9rI1BreefYI3H0qpAQ0PCnwakRb1xH0Z39xtfpDv7kdmaBFh
Xec3ps21UynUhLrSGHILL21Tk2cLaX96gpO4+yP3hHgiCCSjE0OkS3wq0DwDTQ6Ae3dtw6iYHV3O
Vuc7K3bAyOuMZWr0LWn4hQal78rpbuZwi0gxIloV1dsYXZdDcUI1SZCCsU1ho3ak+5JokGKqql4z
8mmEOxRRmKt7l1P7pwiebUXe32WAJk98EXfZzoHajeMh4PioMaZHuwi+ZEzBHs9dGKwB8RbV+VY0
GXWPSLeL570bUB85FgjO3HbqFYCv4/iFXdzR2JzJlp8OkWDXlmOv6VbBpc/InGqPKH8WbjGZO5f8
euMO/ClXCtLDR7lASkoLFTCZHk5/9M8Uc4IvI0XzJ/r6ihhV55obu6UxRhy39xqeZt8gpM6SIsOX
ALofHezu7hk1ijZ2Gjj3zhLIjHS/2/k5/6LZC7dBeNfnX0P9/RF6CL7JfIe8d5Fl/FuS87aH84G3
X/4vRLjoWpZ1Q/LommZOhfX4C2GJwqznwIx7+uu+nj14XvYUjMSbv5WLGQxpO7+JezeORyW2zkGL
0SgNWLZr5kRLTEmSF1NKt2fj4tiBSLUMb5M47m/y+nE2n9hTWn6o2WhXfXy1hYGJpGZsrGV5xmxc
FNpc+/B6BrYF8YQIdZwF0yrObrQWBwHwkI8edFS3KuHsFgJ4BW0OKnRZA5PqKqoG0oRgH/fN0umb
AL1dGKuc+288fSuUZavyPOtGQ3/u6yKklw0HTeNRFP0mkt9NUU2Pr+syjBQe7pjeEfu6SDp5mZEF
6yqUgaboFIKuM9tKIWyd2Gbrf5brAMdX5/Yg/r7O4nM2PtbudnLpeCkFSQIWQv80HwG6JADQ1ymp
OUgw6SmPD6JRIoOl+Y1YwX2gFOzphCsXjheDeqJoIAFTEiq67nFBrUCmbodzUT3DPX5ja1lOhMrG
vLz7kCDzydPhMqpBWO0XE6O9yceBpWosnmxS61sKv2j7V9HxNdsGWClIowd/on2zjNrlLHPvizMe
/u5mnUWG2y00vZBQCFevmqpeCHzMFdWq/9hnD9++KSd1eRMn82Irnw3j53NpbZ+ghpYyLZQEmsOy
UlROheKDAgO6APgvQcxLVJOImDxFSqPvuDsVCd2t3neIRI/FTTbGlX4/PDmxQAtmS1+kL/7wiLGK
rMQkYqdIJDFXSBZOd57bfi8VEGxQhgS3RDiS7YEYy7RI35F8zvC2MRhkeN8UMVicq2ZYTtt7XZS+
8OUwSBLL1MeZE18ElRruitnjg7nzZ/+JvsOu15Y+tU/CwGHdWD2LoNjdy71ox0zoLKMOumKurYM/
BAWZ3jwF6WIdINKM+muJp5om9kmhRaOy20XlqJLdf7iCKxHBLmqMABuF2NrvDYsFTuQDaXamumj1
PkPAOwZsl0Q/9nDXAEyYilT7m0OvCJahqaJsSSNMtd8lGj5niLzJ6gvbrgaMpEBrC6OFdbhAYKaY
Vi2omU1xkIrwosGjctAAMPX7UuetCEWlUoLYIzjHJQ/8bBc4LAwr4Me6qNpoyM1pidYpi3dmIzgQ
F4cBSIfJuNTaj8ZpVBfANcvCURIafErzt4nWLhARiC6GK93/jbRPNHWE6obGO/3m/hm5yo+uWLlb
4AjiqQh5Va2vZT8ZAymRg9JdaI1hXWFtTgURrK+U9UqDtlQY5GEBFwk+lkiL0/HvISyjsXDqm57D
TFgrG2nHXbNeecTHsu6azZ4UgHHlaV7qO9dWrEM+FvfmLbsyT9o+DYkqcLtKG3S/MBza4IGUujhf
eSxVs1RUUUJx5ag+KV5dvCLG7z/jK5NVIbH1FY1Xeko2da+K14mRCDekuhHkk6z3Kq/z6Q8/BBWs
O5IWoyx5liRQV6E0nQaPczSyN+LSXrkaUqy8N78+RYN64C9Z7ifIl8OrpGjVjTrEXIo3fnahxEZR
HK47YNpeo3h8iPebK/fC5BnfpnL+tB/b/odqcC8K2L1jERyta/eaVi8iv4qkH9UJ78oPbmHy/uME
xu1IT0H7x+5tOuYphsVmuV3tKjzOVK1eTZt2Cj1N8VKNFpQWR6IVda2Cmv73pwrakcHRBJnZtEOK
6WUBlLl0rogInKEMLy1xiXrAmAQI7qHBe9fJJqdzCFPK2d62gr05iC1EV0y5EGoJIPBC4qxr/ul1
KlCCi3R2NOIjA9B8zl3NNwuWUAR9WwB3xFr5QfRMn5gOYNYoL7LsS9titfGKSWQVqRszrhVp7mD+
nUz8ibF+zEdPH4l1Md8UZw6m7UiLgTxPqEGxPxeywmacoqGWf0qNF4Rsc2SpTrpXGjuE9zGe0lLw
hkcGeIzUaojaTzRJRX+tKreUEVPxFvIgzb0kxWT6VN+l67XQYldRZ5KtFiKPrh9w0imBjQ635TDk
nLq3J0dt/b6KHUgpTVi0FUs+25K7hcyNnFoXGmeRy0U6fMcdJathA3FYu1BG9U7L5pjSQVo8ZspO
xMTzuw0Z3NoHAxzQyi5I9wUsLrTfblRSkTB/l27/izgzv5DeYyuoDUFzAk+KUnv+fnwqCLud8kjn
ZWcGewwmzGQEOsMEduGVB+0KhMT3MeHLS+91L3amdAA8YDeZj9/e55CA8SXHRao1AFxuukoHa/r7
MOaNzDiPtjAj1z1enrx2uppl1qJQJxKCSJL/6g+gmTc46oyN4g5GfCOv1WJCXeio9HHLdbetKtBh
kzY/R223fPjwWrrHXoYiSnwHR9Te1XKRE9kOx+IvJljcHSlHhC5vUj86PPnqTruLTBN27JjAly0c
MU2oc2MF3vwxanlDc+H2GZ9TjxOzzKiLodo1+Jtyw+qH1QoFPvn1P+KkWonK8J8gse7VzVcKcqFh
d1eZ5iFqClMOwec3T1T6+awHDepJfjDgNEJfdN3LNrz5dAVIpFi1lFdL77zMiA2+B49mj31a+HzC
cItPlBzGENDEO/9i1HfeHfVY8ozLko/kP628xALwM0JbFTiDANLgTqHVjmuyI95sslYhR4hQDKX3
tFruTQDLsXyjNlqQGYg/LaQCv2yDmdhGtMRYl6PC+U6S91uspJFgfWiFmyb7oDKyJHa8dyjjbx9E
cH7ewNaHEQ5xir4cFp7jIY6poGIk6HQV3t2uMcGkbihxd1EixJhlLWU8aA0Fp0p9PL2SHkWkUIms
c3SXThPW8ejs/Row5iudJkgVwJtt6TtqB97zAn0SzPhMMZ6sVGWQpGDM324sasRZJVBc+VZI2g1J
fodr96aijHvqP2KE7csRsBRzBVyIcBt83vl2YGydeXQhZD41a68WgNHHkw5ZLE/ih65SyaKak5XA
s6dezSeYwzhD3l3JHQ8k0ZNk4UrFq3nGIfEkoYGiUjPK9d+GDbDx+3U5NzCjn89NqlpQFBduVs7K
Q+WTXR8IDeAt2lZJ1Hj1eF0B4KfRs7UytrPcuZ3WnJH9PZjwrPNyNvOozvVWG2qPZQehxwrgy//c
wJoHrg/dwbiXBIhKBWDwb57TwMj2wRnNN2qWVdQB1E62xgb4F7OXvv8J3JbFQxIjuGGS8Stt5DfF
spZ9ynCNw48ag7VWRhLt5eOjtUIelo1DfgrrogjHlrcRflVZzJX6CFYD4tbOAKJJEHQZEwlUmJQO
fmuMmr5CJ64K55rU49XWHv2NplLxNbtPMM72TwzL25FNuSoHjNjII8qjhC7DtIoCNfd/bhOk5r7r
b5gagLnyxSxnspFktSgVSQDTFVO+doCbrO7zq0jh3vRDBNPJBd5Jh4zQgYs5KH+MB2NrZqSoJsOm
vcdnxJ0hq2gKW4j7zjS3Zud1YZ9ltU5U7181L3I2/KmbOLdXviIjn938i094MyDHRibG/UT7WQtw
kiO4hLB4iT5dmLvW3BQyaoiJf6e81MKukdS7l6KITRYNYXmspMkZm0O+Rg3y9W4UtFxr2y/SCazF
89Atcfu17U8Vyy8cI1ORhbFJVWDxKge0Ik72w00R2wtNLOQKyRVpaUjAv2jl8bDjiKPevIz1O/Q5
m6QNi3xb5sVXROfZfZpbShMk6yviZFSgwUWmNDA5oJJTBHsfZG94rtNmW+Id6HyGTYYCQnlf6ca1
VC405lhLx32joIpbI++kCOe5PVHfAKlBV2b/o8iOnGsqVl1YmDwSjTdBPYEuuhOVatln3lDK0riH
P/ZfXR489V/jqDx6tTDj0NIWUWtJSxwNVLGoYNxEXK+1OYWINZYQNh8BHBIvAT8F5oiM6K+Et/Qg
csTsWo8uVs9kXlvA1i83otaUdQTsrNNPuN4UXcefuRvuJoPuZR3b/c+kGkr0EJm7lyqTSMUgRgpE
xH8Gd/tzYeenxdO5N5LWk1zGjeRP3HgxjGE9hytsn1lQ/B0hbFXeeFTITFRvkNZPegbmV0PusdZJ
3uVsfJRTIlT0xRhEJdATGcs0/3Ey/5+7ZUvBef/7uy3LR/waqQLggpTro6cIAH7y/T4m+UPSqQJ1
4OrVy2/Z/EVY/BarFz4ZkxvzlWm77xYz+TVhNRXIUzP1JM53xIjyyxg9F6M4CAv48BM4oFy1FkfO
ORSlCwIuW5CGELjNfzxwvD12EC7EoFMfGWkUHHfNFl7ZFBvQX1vUJANFWZCUYcf+J1B7MkH8ndl2
ij9NEDu4UKBYFxP5n7bhRtUVXhz+wgbJ6DadQM+ImKUl/gpTCzorsnfMSph6ApaOkdNlh5kRW7xU
oOw6vK3l4sr2BEggpiGexH9PUIOpb64EuPXlo00+sOhmpSGiSwBtXcJWaUMAiOdGiYp29in524m3
cI5gHL8EGxkUeMiDGBSEKwgBM3awV5VDiJZZOiSdPN3Vyz2bqo25uaKWfq1ibSejPcw+zQk3TTaD
bRK66GMgCEuX0u6OiO9X8DtnWv623cPE5t4HZJPAF5WTCIgtuTiC9ZLDpo/J+zNmcmQDbfq+9Pvt
2Ap+6zsYo6CHezggZwUhLub8kpDLAP43ec9f4VQ93Kl7ubtjFwGyEx8XUTSaT0eIxV+bz2Fy5zTm
R+Zu/ZVPvxfGoL1OUaJxVPfRbSKOLr6humT+6usIDJjrjsrJKNEAtKLpY4dB5Xa3xaO1C4Qawivh
ibxl9yCSEKSIVuO2CDXsaTt7iPxI+OkmoNwUKW7QLj5FF5BR3pTJ4i8v8fkIkXLnU75yc+/nHjPN
6GrkcvJr2671vXWZ6Wi7wQnoYFkkqNEP+YfAAHaZrnUn3Io5Tp5pXbih3Tw7fEFCzAAZITi4J7JI
DTqikeieJfbutFrB7BKIiU8NZA5G4otYZ9wqOD3vchKL2TELP1TQ7VGv0qIJcF6SCirUUxP7+KlJ
iOsb9iM/1cLclogYM3FoqzNa9LFN+s5K9na3kCUQovogSWmfw4kjWr0sG9mPLfyYrc1+74nBGoXK
cftYL2EhtjAcYIIOd4GO9T4vn3yzl8iErZ83Y8DuHeq1t3CtB6le8j3io/z8jyC6IAuEejvyeSYB
Kl1OCZc/XzVmS9trErjk9E8YWFXmZGfYgkTCHxnQXMOnq27YhLYlwnSpwAT5+de1Comzbc4dfG7k
Av5rthUscP3oVg7MGVKgBs4Wlf+Wm7YLV8ZP3shKW0p36wI1Lwu4OASWEaj2f8BE1FmPfxQZIfzj
wCBrXN2Qa/m7J1DamSq7cbe8SZEn/qZQAqBK8at0K1sJptqGFZpynGJ54hvlx6yYVigAhGPfOP3y
5Xv5spLTDXVkqtCQbw+5OkAGByg2UhCkULjptwS2yjE/WxcEh9wLL48Vi1+86zM0Tx4ABWXnBUDw
5pheRFgIHSP/EwFtKHjdj3j5uy23P7wrL0DcQ+AugLBUWgOW3gRDJ5SIvWE/EEgIDFqE66kyJu/y
QD1DzYfvUZ5aPkgLi26rbDyxGcMcKEdoxrWTzo9V2SFTA2a19fB3akwirNGFQzJoRoCkVhcq5PD2
aWDpyep58NtU4S1fEPJD0gpqYi571zV+qPu00uuuZmYj86N0KqMPO8vZTIhabvtR8sODY5aDHOUM
nRfxFNGgNIJVafsgNAoS15R/RikYY2p4M/jwt4NvStY++yXvqxws4iHgeVe7ko/E8PI73Z+LyPfO
u63VQVl1yzxs7x2ZmMlpHzH9m8BC3+ZXauaBt+AvJTUKSHgwX8b/h/lmRuOgbxKCdkSUawFY0y+A
+pt91+PqX6aIHK9r2k74MJ6vxJGT8rvFSWitY56cTfR3k7v86oIDOIQ6WG+PenxUNhS7Y+5KLBFq
5lqG3qC9ynbo8a9Cd3nnN4ApfYSAE/KHhPlr0mlbl6ojdXupesGYQDjQ5PHfq5THXxXUzOhd/OLZ
XICZEnARvGIRtqYd8N4LU00rqIBvOOB8uiV52IIo7Zyn1Mwz4V62ZnhrwjgD4Sl16aWVmC/255LS
Cxk4zXoTp1i/73wvSXKVOhVAFKab8n6fMD3mtM1Kfv9PKA2CCBCTw+/oglwoTAqa2V/9hE+hxb7K
Md7b1BYKunDIyVRibFJyUU8iNeEEUQZ0rKwE8IuOMqfMz99RVaUqVHmtTwHZYIIAvdSX+uR71I2E
tp6ZEKpS3un/Hm1Bh0hLO/YuTBMswtRT/lrpWft5j/hSATLLNz6l0mvx40tGcPgrJjSWMJt/p2H9
4LxlGc0TUo0AtBtKqb8HiHdvhr3DsyAn5RVCoKoOyKJbYlffgQTYiJ0DUf1ml64xf+mtojYe6pjg
I8uX3W3CkraLOl9KTCIEPPvUpsKqbfwSW7djPOespH5qCHcWMhXsNr9zkF0oxzialHDv+3RN2PuJ
z+5Bl4OySh9h4kS/9mhycJwfqSsyHce/tqXcr1QwZU57/E8hgI6YEknUQJQaG1jSXTLVYPCNY22P
uRlF1wOQKgzbB5JBFrZdhW0lp7sxiFJtCnyb27+F3pVO3RSHg88Z02rrQUVLK6U4myo4Tl7vhOCt
FCS2w7e0ypzOg6oWXHC2MR8O/Io8GGnZim3HFnN/3IbzuiwRBwQfcuX/PnJPC88FYY74ZsyNIe79
rb/L/gISU4lF2BJZMlBoiBcmnObFSedupu5jPfIyTq7R0/SQOH3WLz/mK0pzqgtkQWptxd3VoDC4
1oRo+zmpIOgqEH+uIEyJY1SWN5XCid57D2U5dijeRAzCb2xD6eCG6jPzDqwPmtUxpzYMa0oEG9lv
kdqCvB1teG7WPrw+4101+TlPT3RU68/o0Um22EPamL1WnrrL8MnZlxTl0Gxw65kgR+jv1w3gyjmj
WJ9p1150FlkW9mSWtabLBa1kdmZQuXoiELu5gAssrJY50XMX0wXpvpZQlmTeL8Rp+Odm/l/xP+Rq
I1WK23C/dr86k9gw8AfItZ/xLSHM8OAotOCPWutCxr1i87fNJEhRYWqVYyiQ9PsDsnnQ/7hMFNvI
M4ddRg+DvubGsy3aoTCJFCYppLRd9noCDuwotcmQ4JIyTAxo1BAEFURvXksWguHh1QDOxkxBWCcm
qOJHDOCyukRmcwsDcRAveM69ZHgAePZJbwN7LRyM9sHkpS8DmCk7ZJSbOF9Ra9rlNImhE3mGZTpc
8TE7c793w2qFsr1RdBhG0VtHoI0dPkF2KMp5aPAt/hU/46nChd9/ofk0qDdQtqOQ8RDYp092r53M
PpIRQk2noK9CtkxVNHawY3cDf/sXWpCzc1wAn4M9jkpVgoy3cde6WPlI93OuPjEGArwFIV6TXotb
VZR8TuJ3DHGg22msHt6nPCOPJmFE2yqJlmMbJZRJciWjwlzKWL6XQBDpgOZauUVknEAtp7YobRx/
Cfv8L/teAf+Rj9WL32eIkj3CKrGa2Gbb27VhlQcN1CJgM9c//7FCUZBjDrxwHhLmo6j5tZoLcYxw
BST66GiEznfmtTgNd3/Z1W6yr2CcRApLvZKCjfcBjcDJM5Awew6kSlJ6ZjMvqGOIt/wZCQNiERzF
TSPl3hhPhfFQmGO79femIwzZEI+knQDu9f05EQL8IRigmJaxqztQu3Td8aG3dw1ECOmbMryNZsS1
JHYIGmr/4NbO2YZTaSUR/johcGzmzVW5zoIFl0l8RRpml3Ut/wWTAUWNhRZ2lSffDi7X0eSV5+Kd
aOIAriklb2rPj93ClhgJoyVzCxsNf20MxdZd+AiKog4R4UqNhRdnrDmAI874AoiZUWcLKOsNltAT
4GaIeCAw5DMoRbvoFINuXQNTM9ul/9Tn+OL8c7I0fAhG7TXj3Yr2Jtx3+aShG5v8jTa1lYPDJ86o
kclTwhy0NyLttlNsNP7wZtDR6DoSQvCQEZTEwfk7P5MW0KYHgLt8LLMdUIj//fPi4ZA+pWi4DjKF
EUHVc9y5+xXwGjuykyElmSw4Ynq6wM9t8EgNQsp4s/Si6LbnhyxcHxWntzWTYvFBbDIooYHZNn8t
iMrcvIUCysU1vs0u18wku6EIBMDyUMAncslIZELmLn7dr7aIEJjUkrGZPjc0DY5tssKNOHYMNpEr
N0nZNR4A02Qksp5qr+0W6R75uQb+i2bjKBh+EbtKReUl+yd18kvuH2e8X55KxV81Qysf/R6Bfb5w
b4rtDFFRk5qMV/AGaWx1FIsM7cSn3DVp+rlBWpE0le0pLKfD9iXLxfvxPp3A5YahKG1Nm1wR83j2
h56GV0qzV5AeycUmN1UP6gZYN4z/VHb3dgkzGbRVX8IEajsBwVGj252V/zZiyhmdwaW/VSAH99py
f1sXDnDn4LWOyE/68bK6zgV3e+VzOeskeuu6ou9KeW9DuSb3tPWbYiFYKqX3qC4vXBSloKVGQDiY
HzD/5fbDSX4S7J1XyHUqPHbewjJ/jBSuw1A4HzRSffyivmj/xksONbTc/lPtDAdETqI8AVMot5Qf
tIszZ7YCAbrKhXzFrtwKmHEtf7X6jAdmyk6+aKhr5yfEM9kIWWiOkyzRBys5cG5/bcQBxLdcOEaP
xO3Dj/U787U7zKKIoFqo82BBeOHimMaz7Q3IxOt0BkJ9hP3EwGP+w/PjszPfo33eZhJIm2pt73t2
XM8NGqaGmUxiypVKKqQ8briWs9Z0SI5wuiZo8nzgWWMOw17o8yKNLgc+vxwZJBocOpZ9t0EmP56T
By2TBo1wVUZ/oHscbNoJ3HJFtuBG96UF9QGIQ8whjmEZ0VYp6yJVWfNHIV0JlIm+33CO56xbHB99
g7+uhJliZMR6AIfOI1YEo8ECBbS2QsPC20RujaetbZSTxcPr7OGsW6L0ZJrRj3xFhdRVrB5BLOMY
Cq0q7JX8BWQeSb4G8/evmc8CfO7KeeL4oLXjx8mOUokGqb5IxffdTPTTd+ddD8lchXH/3GpMP/2D
67XbJbaJc2OrbsNSUxIayj8pWaAzm2cmC53ArSPXjnOxlE6b+84kA879ZyZe5gpE0C+n8HQ47yEh
45zFRDUOuttecRt+0vD2A/ZTSqUqPrNfs1SqLsfDOOPd/TOKPOwvtmmXzqdS+NvYE8Z99yGBecfI
izp7N+YaTvEKR9swmNQskOjeh5l0+XSq1lQNAq86dSFo/lJOZV7ds+KuUPjLuumZwgAD14XplB6f
XYxjZSM2kMQTQnm1phRT/7bEtZ9HDHGIvRmxoLUHd3aLWv/UnyUJupJY6JZFk10QtLhu0ERIqJ83
iHHRTpJJbcKBvhkdvmNh7MAN6+8yWYPQLV40ZPY4IBz1kZBopQkBglLrsylbRUd3dgSmkGbUtUTl
IPTVcHEfikIdVAOjo5jmU56EEC3PhG9l9ZZ6q/CbmQP5LwD/uwapz1b34DWiXa2CxLV6W2QWZrkv
dJ8dQo73cgOBQdt+M0vdYu0+d86BQO/QdvVBZt6MwGNHShBeaB0HLGKBG/ohAOMVtjCo+IGetean
1lyTWLFOVfpOw333rAVESvijUftiC+ZNSYdpwdTMk9wAInz4tkJGw/umDHqqzO2BQ+As39ZVBJQ4
1GkBO54tGbHAa831MUkckxozitPxqbXvcdpr7k/1WZxMAwTOmlksahEnZNLVhh99MZ0qx/kveOKe
VMOwAF7+pVgvkOu8bxa767EvXxRBkVdFW9J+G4KBWUtj+rO//oPJ4A2QIdb8qx8uKoTRrfbmmSdk
bbTPOZTP5s34YeM0KHsVd7263Sk4Y1qBcC8eY+KnhjatkTyBwc07CpPyVYlIRG/9HtXrg/ClrSQ0
BiLuX/HXWwYAWj4rAecGitd2YGWhILi6UOJlb4biaQyxxG36JYkp6P4HIFHajWBMmka7g4Q+i6c8
dFkRlJjMuehle8wTEg5C3vVYcr8+yV/yrGkLB6gFr1w3kXGjsc4r0dgzxf7985Rk6XEKoN3QMDBK
EGW7EThNfGdsLBe1SfMSah/gjdt6zJlfF1hMuVZqMfhgxDB8n0GANcvJaoqpnQp18EqLE7hEn6P0
JQgG0qMEyAacUKkqwwlTDOn2T8fQFO9YnM+DgZ1uXkQf+yFVsLODygM18pTHeLzzQkC5y4Knmo0b
9EoJnLssoaK7Y4O+KRrxnppXeMxrWztMYfa1ehrd5wwtnA67V47nRscxq6Y4tk4imD6xP4q/zLuf
1bdwSPPCsA4U/uevE+6HOMOjAYan90fkBaFfwWV46iE68QV+D8LZAknEsJTr4Lw2NFQl1Kv3CIgj
FH7PBX7vaBSECzKT9FlMa1f0J2DdOAhdgUWPY6dExD0rT6sm6JpTvUODMXb2vdpY0urFEppnAUd1
4QHRE2VJeIAkio2YXTn8uhwg1M4S9POzJgcVz/ytGWAO2S3P7bjyUvjaCYPglNr1d02U2cFqDHQ7
aKvvBx50VSYxfYRmzA0m+JMql6Ij3kPQ6a+embHPHcRiAlgNqSKOfw9fnV6XiyXonG0Td249dek7
mB1uNbFRAz+IpM8TGczvkp9m0jANyhxQwSr5d1SLp+5ZA9XjfNvXiqFW6l5VLZw26grtwvOrB2+V
OaDPD2p1KKxZY2NAQEhSii8mdnfFcGbz6PW0+xDlk6Q0qc9EV0kwZ/56fO6VeRPavbihcQ4+zRuH
NfA4dX2RvWZ/WC9/Iiul58bmvyw0Pc8hA6jNEzcm28aqSIhWjzi19cLxvYNH5v5Rv5YEjQ/Tm6PJ
OPgINJhwNN/y1pC7T0g34bV+QcQmWABN+N2c0u9F6u4HUWkJ2E867IB2tuur5rT3QnRIBH59yyUZ
UfxuQgyMVKv8ToYb8YiVlgttO6k6IjFifZiEoBGyEjqvTECkTduwlEdKcJdsfGHkM+BQht+sVexD
IHkCtOg7zNpTmw2nAP0WmXqh5iO2266iT4XE/evAWgnQ/2iTEuf8uSBQ8+9JiW0dH+RPVnkpFSQh
k087smxMVhVoLKkzmVcap5G/RnJmC8ZXu452kKiVC9xQ0Aef2xl7lF2SDTxsIc8lIpdJYlsDMmZ8
BSr0waPxQJINFqcsFwWM0WPw9/NBfpSQIoFRvsgmly2mA2T+tzmHIYW6k9fYe2ZCmGJhVStFy+lR
ppToQgNXqzIu7qdG+aNbtD0XCu0GpwI7x+mwNyahH5b1zAqenD9giMN8EVlqlFKJbPPkPjE3tTcB
8GWrgaJxTRVcwegD7R+ZYd3hUxQICzeaTQkBiwhBuLupWpNhWM9OQ3BNlLscDj/1Y2YJpml3hzsI
BZBHULA6mgiVRvDs8zZ146i96QOxCk5/RvjoKqhIY/lvxeXIvtLyiGE4a2bUKYNiBvWeVQXrH0I9
TS07f/8eILCmsupxmWGer6/6CBsYjiJKHoRA4wJhIJ3fr5ataA3qmn048r7+zUuiWaOYI+ZGp7hM
url8jz2O132vM79ZOgZ3IXg+fL0rdJduqTsoNRmJYv1SkZrIVAgMQUMv10RBkJnhPDqclbErRPjK
ChfgOnTjYsHh3poLQM/iNNoyzIaLyQAvtIsU3QNjkzNaBDcmDauw04WGDy93BChR+ToEgtnoAVSx
JPFAA1ljEGkyl1+pKRjPoD16sHvhwq3XnmnhX5rI/eXL+MozccjYY2+g950pfv2ZOl6W+vrfhDDF
HqzfwlWm4TzylIn7WPDWMVJNyAJZrPiDMstbyPukxyaIzkfDB/MDWOEldaGqpmU7Y2TbxTpYWcOg
AblZsFbptFy0nTuLyFbDXoeS0yBPTK5tukmSf4vcGxtno62C37XBwNmlA6OmRbcglGFvlU5iEzQy
IlR0tja3YEiTr0bDLBArdBIWEYfqdSS1Sy3WYHipVotwPY1Z5j2/YwRrIF2UE1cVwEwcmCfNmqKY
PuLt5Oo6FNJ4mdgkA+aGJX9KBkDJxb2xLyTfjXpLt1lz0R0XU/JYy1jJP1YtMiIqknETcXQjop/E
lqH10i9XxtLcJMPCmMvE96XaNPEe3ozlozTDYbBRw7lALJU/HqStE4s93I3KMgwZbKC5tuQDMiOk
MeX04to/lrSTkymJdjGWHZCp3vCYHGnLCN1B4rwEKpU5x7wSBYtq8+wWi5FUottLew5kdvli57P7
lx1L5+UBlwoui3+ocYgpLKQRjHwUmSgEBffaPKxrQvjeFHe/ZRqIA83kogmoOXSh1sMtwsVMuEfY
KRWNirAQN4S1vvF2sajqPE1ocDAHy1SuNuTLWXdH6Krq80D5lPQTaGFDRjNnYb05n8o0c20KZNLe
Y1MVWLBlqfwqdEAawP+sOMRMABOEpFEG7eFxVhYmBt7a6U8iyNbR/v+NVjmMln040SeYHrzqGiuT
EVaZLokxIgh0+VmibDdYO5qWWDwMRjLzxchqcxgH/IpUNxX58hI/VOCEzCMQwaSkJEfvZOBgOYeF
DSYCMJAh+6B8ih6DIco+uY0nTwATlXK6XB6athArD4fooyeq09vomFfI8BTVMsu75D1O2a0OLp11
ZkdNiIWW9AzKKNUKG1iEPI6yFgBa8c1RGOMq4bby6LI17toT7dDF+gGX+POOJ0mtYr5pp49uUGIe
fDqfvatP7u6NFm17LY/On2rz5yi+9L0shBxhKHfiQFFwmzbmGxyVOEntZGklhuP6LxvwSF3/g0Xw
DqL19kaUWxsP2rWJRfhwJ5HOS9LP43PnOAs/aaDiot4m2Ckzz5cdVFvTdidmQZ0QvRHVhqTaJHfO
Y2GKrRyE+/AMyP4CkLsyoLp1fdWzT0vHk2RhSp5JEqur0U3sZ6kkzi2eet8HsOWX2uFgFWLkJ1mF
9h102HxR403bRgnYJOihIqmSr60QNzbLBOE3sRc9eO00M3GFtuTWy7xiHnzIAX8tuztUck8CoxdE
8kjwiVbmrHqWTfnhR/3TBgUYUp38vZ3lIMV8++2L8nMyafJ/PL1xTc/M7vkXtOsx3SPbtm/4sAqI
ntFpSa1Wae+lcjBMBZnOhiiqiD+Ukr6Ywi8z+QjN7ewpAzIBp4mEzGzuDa9YLbeYVnsi5u5fzFJg
G8ay+iKYsSK603QXLeHTD759OmGhMqT9KK3LcpBTLEIAKpkuSUsdsQvvlDLFNrMD5HI11zKa62aI
ERv2Kt273sKH2XZugW0TfPvKDVZfN0JVcf5E5GNe3HONjM37DMML3IUHDdVh1+751KLOJ7V6VT5n
eMeKkKNRO+rWhRY714T2rodoagTbyfeCQKC9Cu8k4KjOHPkqWEQ7n1tRCkzgXPykfY7b1q2tg4ng
xQWqSPcVWMNnQAfTR6lsYkbw5NK5dUgjYsBeycbPf6FMfeVDpeEg/ZBxAat23HH84aEqlSSo276s
e9Eus9LXxI8Tg+H28es/oqxH7b0iry2MmBLdlnpgo9bj1pHQES7wWMKBOIrmotZN5L3DGv2lR8WN
2kJZK0ZbADvNaLz67GsRjkzqgrZEP0QJxpF/V7Sv5S6OKbtBtIOATB2QOnCZ8E8bZUNkGlEyS8nN
RvhDjVdrxd/xg2NfVjW+l42bmxtAxN6AgzkVQ1Gly3xXkAyh/Y8R9AUzygLE6nqyY5p4PSyDAWmy
w7ukDEHh/rZafdveVbWzrpjZpNcct2lYPKlGBcID+eSQ3T30ukOF7W3aFkH3K/wY807gD2zn9moc
rs2XRxL6mguH3T1ejOEbFmpDXQ8MY2pvEDgKm1pZnVFg4vgbJb1uyv+3PdyiiLO0ZriyowLfCdNV
fm1WHz4Q53cJY8Bx/GXKsTJ9zEzyMTi+Hnz+/cDa5W7Z2lswv8QhIteTDmw6SrbROjlZU3oJ91VR
QZbruXFA5fzqkLRo0AumxN6AV1L3pRmN7sTDbbZ7jirmL30gM+XJyoOnR54uWysLpxOpwpT3vUYP
YVIqoIOtyoFqA7gQRw3EBOqm30TmOEn9aOZJzjElzfcTlQdD6QnCBLSjGlwu0Siwa4nOCteWNca7
yo7J1pTrCx5zoP4aLSVUgeTmkmucUmjWvBOxjqUFxpLzBu3X3aiKRtZPhrLHTdmd0EK1UVdul/TP
4ItXIxpIvm5oA4/kBtbt/WIu4Wf6L+/FtqN2S26nNubR8Ay5on54H6H9fGxL72WSOUN26wcCD7qK
BK9V/Q5qiM0Mx6CZ9UB+rf9oIL61UR6Hh3FCJzQA6Vt2SX7J5DTbabyWcUEsY3UZ+NO/VbFIJ8hv
1UCJ6cbWjiux/Ln6KIvAP0gdRWNbp3jzRXz2eiQEmcmyyIHDgd1y1H/NnsbTQhrsGURgoZCncb8Y
sFqsrMqXohL12P04rlcPo9UghyrO+585PbIk8RYb1V9fVhB8g4QuGe07KjK9L8qJUk9/xDzyZMh2
bV5tm+J+SIlWlY+BRhnDY3rU8mrqWt/vVI6v1NWV67znBkOssBJ9iLDmu4TvRlIgClTEAEVP3cn1
Dqv8OwfMZrtALg3ydjw2XYIr3d8GCjc52M6nqiXhq9jV70HGjJ9YxJYxxLcZkoJ9hNMGc1Xo53QQ
uJMOFWOe+xiPm633AcVkagCrFoZnzl2RHBN79n26V9MMp6djyPJhHt4t0WBdLbCZUR0Ka7pQulQI
JD32O0CUGfKMCa9+V8K2dEX2DAD4AZuPMNDKo/XMO4rAlySshmAyfquJijHSImFxdM2AP1fK36J5
5TOVDEvQW08NCv1syaOqNtggL0lDKE/RkW76Hbsm82Jeqv2knFTBgy7thb0UwjaxVqKYWFI2nKgY
B8Yu1B1+Dxm5l7SzcIo42uwfmOAr/qa3FsZ6WAU2chosvgm9+Vj2tY1o7hWYn6v3liNxIsiPzzNR
mgAjSpwJnepfey5Vol26Tu+91ryLMh6JF6XxkiXyGYgwTgPFlmtSzNDglK8qlddlFMrdtZKlONqa
VKc2QtniKDx26Yt8qWaQRA6m+ccLRs/JzNkcDoWZd3ibWQnc/XBCbL1GwavXPsPrmHMk7Clj+PcN
22NR8LHNbduGGTlTqXyGDQKLQ3MdHX+H09CaeJsOXGnVCZxyh9LqGNEgVrGAItn5LR2LzC1ULZst
Bxo4K4JSN6YZ1HZ37TUVwyW7H3sfurJJZRYIIOFlPEazrlG97dsqyjIsPF+MZPqWAJOkDNw7fBE8
JBCMZmpUXABe8DGeCx/YGmDFzDaADvXarTzHDTsV1HkoIqj6F5k4AvuUncRKNJTl2Q9FD/KhIvao
LWMBYvfTPWiawrd/Uv6h9W/lPxOkIq7RARFH2kREdcbq8nr+4yFaxoMYaTvWYIlbWQA6qikwmJFy
FK94pKLYjz2HaF+W4WXVvx8Jr08+qEt0sJWCjwHUKK4dQ/9dzHHprYGqCGw0CCZeFY4laAr1SKsw
lfjuGJ/Oup0ZxmbdrU1L0YssXWRh4TvjIdP8xn8SdV74+vbyOV5M3OJX7zbUlD642DS//cYDjF1w
C66HgE9E3145TRnlHSOjq6IC+vvUQGXsTqDJbG6QNTmbvdYQszRA6U2GGdutHG/4Mrbq50/OoRyO
g6XRIyRQVH/Gtf+jOnU1x4sVNHKtJ5mDKVIe2efd08AvD8sFKJ5MjPfDkzRnCfMZ+q1w11ELO2th
CtI19/jonvjKJKmJ0Kq1gQ6mzZLUfCYOt/eotLWkWCxAuKEyCmDaykONvuJefG6AGgl/ODxz61lS
zdA48XXltVC5ORDftkOkerQwh2mp+XafHEFuEeXgPTbKK1leUiVIFQ5ddxJ2A7KWjdp2vgNPoDDz
pMvfqDTCg5L23xesqqo3SZ+4GIrBeccsweNkCTo5aPGN6t4YVPZTeYGVTguK2oBJC7quvgFeWwe3
IW9kZHIjOiJT9wQ4QuPzB31sQ40MoikzMBnMrv8Bn+3E48nUdE9wt7Z4qH15jYX/szCw1NRxZAvG
r+I0GGW6xRK1WJuWAmAxlmGyASX2s2mgquCv7LCOwbunfLAklp1YF+aQ3BstTKwwITP5jI/u9Lvd
v/1PoooSOpIYUML6FnfP22h9zt/d5xrbB/UbAYvVECWRrXFzKvxcSk0Y9xNd39xBpBpNo4EaA3r7
PphwYQ7LDY2W0WC94T0ln5ZfRRgYVwwd3IeG6LJdLgNxF9VYSUc1vMriTyq+WOMxhLoJa3KlqGcN
0Xl1gNjvZ2ghRG3pohcdrQjmR09cA1vfkAZaUqTR5RdJ1CaK4TEcnLYy/Tsy561b5TzE0nrnf6gw
uY3Zj06FXwpPxD2zukhpXym0cIxroCP/mqoTpiD28k/Kc0vIiT2QRZagy+HGMNz4vAqY4hOsplfU
WWjD5E30WkacBa4z4DaUwe0VR7DJFnICWa9ToMAG5mcaonGMkBBiUMW2dOC9V5mDQJG0I2iVWWbw
0A7eCK5bXVS0wXv8yM0m7irHdTP1oZrm4PST7yaataMOg33crH36cAEpmpMMaERIv7gIRXAsYGKt
Vn3+0PHw0PweqxZU8FnDM19gfCTMFfSH7yWDywOYZHS9qeaFtkgSUa8wMZ0j7d3jVaJZzrDFTM0J
I62ZtB+qDDQBUilAGKJJFrUMtr/CDb02uQbWAz7W+Q8s0BThXw2B1vx87Uuey1h6Qi2A8YdRHb0n
X5om8Id1HcjSTnOQm2iu66qzbbjE84ROIqC0ZUK9PIaB7AXAeOKwjUrrakikVcbftoWhexx7tTNW
KMeg7A6ZHHrJjSKaN6lvQtdYkV8U+qS2nLYHA74LTNjflNnoSJJSy2TZUPnvav2WiwCANx9dzJ2a
1Y4ZL8OXoKmysZhJedOvn+f8XZ9U1E3l3SO/5NQo5/KMIU1dpwunVu04d+sTdEuSdvySLBcurIlh
a3UdxXbvP12A5aU5TbSzb6SgMZwH9EWUi/t7vDSSXYem/2nPYnG0JwHMupv5HVxC2Ga0o/YG2Efu
ktZMoTgS5Vwfh5iM3Lf3TA0wT4Q4w81or1OMk5dNsMAWU+avT4/gc4el4yv3sbangWtdRbtMR8zX
DqkScDjDD0+GzRN28DAlM3bUGpVQbRguaLCA+SbK7bOPkPMUkjRpQ2eE6sW4GjUb103tPcYAgAA1
gFnq1DFpz+V/P4YfJY74ypfclN/C/nlOUKedEhsB89+SgQq49k7PC2ozZmBV0oU0+3qcQIyc+Fad
6cxCsJBeMT0jbK9e1+W0qz1VQQHIoY7Aybh8kWSBGwXbUmWXbr1hrMgenN8uqhMQXWZiLU5Diply
xe1JX35qvVYfZajJaED7WH0b6j/7gaqmqtWMYYl+TpZCiQI1bC+khDjWIMcNAdOtqoX6ILxLMVAu
dszN3b1Zl1xDjqEvuUU87919VDH9yQtSoaMtal62OjpVqqPqT4yVtisfSWnIPXsiWOEL7MgkuAEt
t0sXKhG5J/FHPvYQqgTj/B59yhB5T/zc1n4Kt9hkHshwL4ySh8vDcNhQDZ0YiMYScPKsUlk75x5V
WBH3m9Qzug9CX/K1Z5hrKwcC1eq0qMWTdMagVUh4WnWN+jkenYf3ncsJEKHGx5rLBn4tN+O+60ac
jcal83DYr7guRtk5vxzi9AsQ2MP4hdU7nZ6i+pNZpjXb1twp8HKTPZ+YN8uregLvL7xFFu+wZ3G6
jL74jnb9Gdd2pVDykUMs0ni87ILDk4ueELV26rXZbna1NX6gXEpPCx5Sk2r/bzUEw6RqpXzya/p/
n8y11OxGLjSsXT6fpbXTPTnDZD4EArSDD2TGbwZgqintob+V4a+IoAzdTvbiFFDFLMQ6OoOrryZJ
nFicQRBmInYJWRqygutv0Ye/LE6chdmIxE+ZOZT/ELxzm0fGktsejhRWnV8VPfyp7aKYs/jVO9ao
zK2BbCT8dKLtazNRxmPc0krT5W4RDqRuFRKMpRD+FSjCkl+NZXWERva8MWK6Xo006hXorg2vvjgJ
Lg77NQ0VRTpHVhHkuQlxIPw5ADUYsBV2tlwPUeHMyVaq5Wjtn/9bt9a3hpbosJRIQ4dimA55vClh
/4lGpyiJTK0qy6hjph4s04xXq9u0E/UDuHt1wgcWAcc17hpTGSMAXmwyUhNrbRBoBWWMOS4DljUG
ImQ/w0HD16UamD/8JJL49xtPqUFpd530zXY/j3kHq46ZQD4CGg/ptshlS1UDXWN/yzTbYK3xsYN9
WM980irJQFFwo+mzDZhnmUZDlJJNf6iZaZ2GMp3wMJ/SCB7hYDgU6Be8OyNCLSn5GliumsAMReID
EAbb9vITpo3tyUKKAqUyY2ZEZcZ5SU/VBn/m+n+9riZomjEHqvterjZY3SSc2qhNrtT9lSlt+yER
8mvKlEjr+dONxJquIOdIF4BBUZgoMZV6GlGwO8PQphYpFXBOpFQN1PqQL0XKiMY8DRQ5fHVvoFX/
DUpimQlsGOOsJTt1EYuZ0I3k4fgVYa7QSmzP2QYtxiJ+ocLaLipqWMlsdJMKcHsnR2p2uMCFObhy
cXP8opFxreGxfes5gK61GrIjRAG/Loqa4PmWZb2e7Z6+RQ/4gtu4KfKwiCN2gegUaxuW//KKFtds
hueefvQv7b3WCisMv+gX0qgdV8QechPzdda4HD3ySn1ahNnyiGJJPQlWnk8miCOBS0clI5uUseHp
fWlRY743g0Ks4wBQaZqTQypQ9lgU7LxJkKq9yId5lwn5Qqveoniuk5mCMkXs63Si0yqPxZDVhi8v
ZnQYNHK7KPTSEKZRzsWbSR2RGWOJZVMxrnyXsVX/WXr/v9JiTWJK3APowvfIjfsBxvLpmoR0opm5
qR4sS5fd5gDBbBtLpWht4nHyo3JN1egBd+toMG5xoN8aMa06nPejInSEfStmtRsUg82dQUhFRgej
qqnml6b97bFzX2HrTUsuz14spfpI4PJ5Q1lPeYSO4x61xGD2l+KM74lKPVgEjfNyNKgQrVO7gNLD
Bcc5fFb5IKgD7QJf8RVbgYHp8McnxyoElrVv34jblcEI1bzkI7dZnGcZU9rWXIgJzcgN8NydRZ7B
Gl0C367qEz0Hptjkxbh2Tei0KY2Z2BjcpDAzSG+Y7Z28A5pRmYF9ENvWBzRUlNdKV/pRklgnG66Z
L84zIDF7L1hvC5Q1M+THH5bgl6Um+CMW7F5UDEA0XtApKgfz/2pChWiiIYKALrfHpIMDb271T5rQ
ppzKylro/SuAhy7oTvOFyHi3GnA5dZOUuKOeSJSXqiCKLK3Sef3hRDlWNVH9410YQIsFuWFISETb
C3rfok15ps1a1bYrS4A4yaCd6/1gqNo9dppDfF+4FEzQfsWHVjLnS5sTqSuuzfAATVNGeOG13bmG
g5RR3f1fRFcDnJ/3mphpKr7wjI/tJuqoAcflcdZHbSvxKh3KeNa6T676VPJIleBMT1qgf2T1Bwu9
rCVdO625PmubFmhPYc/BoFA7r5j7MEUSa8f/wBxcpTpz/hA5rSNeK2Uq/MtgiYWrjLjJnNwKoIL0
PFyG6h5VNF9WANXqS1Z20YuiwRpCxMRG6sU+92hkO1HmKqtOvHGoQZhUc2vLanqjCf2cL9H6tkA2
A8bOS6pgzvNuRATFc+BNCnKE2yOVyZZ7XWdBzHUK7SxPW6CNUi8acivuE1iUpidx7iB1rBe5jNTA
DuAM8HIYPlPtcnqebLbUjfQePwyZijkQrTWuIOLip1jQgNCydfu9QKj08EP+T6SK+mO3vTIF56uW
c/lU4gtfXtgvgot8HwTB7G7j7b9RmHllyYHyw/Cep7e3mnb5lPsf/8hYf9oO32KwXTjWfnMamASW
N65Vv9hnwcRubSEyrjj7A1N3p8kclF3sKmtdZ5K3gu/S3LA+KmdJ1yKtmxm8yWgIbptp3LxZvFxR
XWdg13Ub3HVih3wAcqbDQ/xeVLEiZ8J0qrx4el0FBQl0BwBlUhsd4yaBGBGGj2xkBudmFedmD6fG
lHgcsSyYc+XaTEqfxJTji/XNISmGUzKIovRyHYJsmphZYbwAL3boXPC2ovTzO6yeoRr2oZhtXr+0
Y+kran1fjSruERxliMX/6CXMxKkssiZ4FFndBwoM163qc58CuOsDbN48ZZ249ZEH3nb08ma6r2Ms
6N5HUgXhXrgNwzKYTBw/fKhn/nw6SKLILu07oJ6HjoK0o/BzZpq/mdc9Nn9IXfY8oICuLNItLuxX
J9TK8lx5wdNDLjpAsTfQ/uEzDxz6N5/r5NfxX4VUCBv10He+OiHIL7v9XsueOGA/KqmJYEN9G3So
5E1wnx69nAXDKSRFyAe52Ws8P6z45wJUKBl9DMtS2Zk05vX9cvG1mZafbapu6RPcb8mRTEBJtsL5
ES66CZxBl7ucwvDIlUUDD9e0nU2GVKBV4ehQoXOqPcaHTRcKVjNicZB6UEzq+P6wAZx0IYMdDi8E
bNWoUL0lgpzzIH1rkyzWdi2VXbP59NoCISn65CWjBaTN9souXlc3n853JrugXMng1GHui5SEXtMS
U2OteVAGk/3IBuWTFfcrvTqzNJCuxEzf/iXN6bhsUB/HDVvswu+GvF2sDhHGtYGLSupLCaFIRtZD
yvV/+Jzig8ZrwGJY7AmeePLReMjZlrSOS5SoZCH+qQqQyoV9eOTrQ1dHUtmKg9ft//tT/Wb2WEGE
sF7ect00WRWib0O41Psq+i1DdyTPaRV6pDccr4BHXxRhGL32ROCVsyUyQOh7FkTVdoRopbvUPmoO
knnSSjpnRECUezBhmO7yYJnx5fymOZQSvKZew7IEVPVAGGZ3D3b1MkJzDqW9Xq//IEwMZHByr/CJ
LxXvodNa9pzvLmfbSfcri4uiv5udA2aKyt3jkGKILknL/ebPvbYuPPZe01/KI33sk+yamwhzqCN0
ECbf9nyR/72I9HZ1CD/WXc2SvfOZbN1KK5vDzfD9ziiK90TQA4lz9fN0CNtE7Dq4fqbzegIJ5ImW
wsWcvZXIqH1KEwnTfiQRzZvx7KibiKae2W+LPfNeIAolJhru3kIFHkj5LgspnI98T0gunowxqdZb
a+ZaSXoHgXPx4M6NbS3hAHxzqjzeHSGaxIQ9FLLt47jVuiT3VZxYhD0qqVagnT2qyURFhuU9E3GT
MrOKFFQzEilcGgZaXf2ekgDUOV0IjtchCEbO/YIt6JCRoTVX52bXYZqOMka9DMLjJxPUDTmbu0E1
M4jkAHO81xTS2zo+1WtvIDqLvrpWdejp1+Au/K2ZWduSjJywKs0Z2y45RMr/5Ts6I0Gcgkzv/Y6A
AmPb3iR1IOLo6tnpwyh6SS8jjkNcg7PIJlQGPewZZKvPYC+fCUrg87Mm1AEG0ZsvwUYwrOj2ID0D
8GDDygk/MBDNyBFtYgeOtGxlmx07qCzwc45OQleY7hBhk1wzF5y5DNQpBctxvvlgs1cygWfumh8f
hxxdc9hfxPM9YjWcRd3YruZy5qrxfUfWrEVR2xj6aFiEIXh00+ME4CmaM1fsCzWju6ROECoqMJL5
f6DlcCwOBmjlOkNdAfVt7QDnTqs7XkJp/wkBzsQ8Il+vwwmEBC377ZxqEfOY0kFHQgPI9rHV2Cqn
9I5K1AYGlghjjH4uttN6fLT4BnKzZF5rpm9P6fU2EH+v0pHDONtFKM6xVbndpcQBpV7qXPkB094Y
W2eTBRl2mKOGgyyXLj25QFTpWD4uSoS8izZe4zZMSSjnyYa0qdqwkvn9tLTym8AqeuUisMIlV4An
Kvf12ScdJF0HKuUGhrczmB0PH3/CVrZNXjCZsXa+eENrtM02d33LpEcqvVownpdS0Tw7dnOV/YMv
kiH+OV6J696CqMGVsJXwaKOacWT+ODpf2rSjQEo8Q+lzev8uRotLPf0R86zEliod4mQaxITPzuDX
VTFHay2rva1yhhiedk0D7bf/Y5e9MnpkLgwK+lCehL2NCbHWoWN0hxi7lgPRdRFYZNkvrUKqw7aL
gMOWWNZ0TmWy4mcF8zZfd81NM4E57z1aZ4TpFHvKaZaE9Fs3ackJT+BOLEDNXQp508NR2bjLrSEt
07jppSWwF+4WDZ0W1IGCl1H/30VSvILgrTNW7+9Wmgr6g4p9gV0HLeEW7Y+tpOxY3RPlJvFAwWca
JH+XF/qXyiXVyGFVd+4qs38hWZhv/O0fnxfKDioHRP3ipg6Qt4KmaT2/zykLr1zMGMZthJjrFrJd
ay204EJEsEmwjbJfy6LmAURLAthb8Ko6gPtDce5JgzYjoUjryFqS94LnOQQ78F9qhqqnoec6Nio1
VuJXZFF0Jc9SJugssl5UlsTWWw1A6F/zfybyPIHBuZ8DzDqluMd3zY1IoPN9VBV0YKEKL/Epak76
Co6b/3rlswqjNFEByvcrW/e1ng2EtWWBFjcH+TP+45geXVB4mIcA4Ub4yxJyU1ZMzc6ueaibjxA2
m3m/t07PfuYVqhWzKw1eKyl62Ur/2X23yGbr986qD1Wv41KvPn5vM5XlLk7/4wAMBsjkfkEPf7bP
d32cMrHp2f9750EuKSzeEfOdrbQz2kceoemDFAmPn0zROcPK6KSr4/tUykxvgy+wDz0a0hdoHlHN
SMs+FC7blv/gp5HpTPP4SUyo0TGB7OOMYSpWlWBcJ7Er8o194wtG7jo7Y6weMPsxyTbWVwgqBDHc
dWdf3oFl/ssfSJldewMdQNzwxRxVgz/d/4cIa8x+C7i2W8qnpQ4DT1s04q2FXxXEIGvJ8yQWU6Zf
b9eqaXx5FN8+tghoZBNzZ3J2w1xe6GESXy1DKKP9XVyUD59rh+XS08ODG+tp51bvFkXxQykcg+cn
LBD6h0vRRuXF8ak+xC9cRSJ8w1bAhFAPvm1cdV72aj2BiFEyPnm+ci3BmYpIVlSM/vnlF34mPNoX
TEF7mEzBJfEwfiMBKQrUXiEWqhxYfvIOd15sOaQdhJjWnrxXLbbAH92DgN+7+w88NQXHfcVW6t26
FIlizr5aKzuOWTkWRACp//g2fnXBykdxcX7ICkk7378joprlOcAwOQ7Pg+0Yycs/uspg/ooXUrHE
BK0yUihY3BQ5xZMyUYMk7WHHvoUSpKxkX/YjXTWEIxPQzC2xkU+zhzpC1g4Hlu2rgL+ApNPu4iib
H7MJUIsPMPhmsKvUSmUxUa0BEtz2FeIeBvTtwHWnL+UAyZFWvrA2DtWEPLENRBmiu7EhIO/pfKlG
PDplpANy6Fp6CVaKKqx66o+sfwcNC97YKMeR5VjiSiU02rB594An1f4yIw9/eJtQtfh2A14FznN0
TsnnrjK02abmuF4uEQbzUezbL6rYBm9BvY+k7YkKYQ02q+NndAiCvzP1+1ucE2foxgIMtTDOa3we
1u2X9Tfab3LjU7+2c+B5Mtz/+elPy5ZtBRnVzPSBcFdKg6uCQ4lv65CsESaqBN+r61zDCoRxZOYI
CtLuKremr4/yZ4p1KsiMcDEnwW2SaR7xHx476JAEkcP4DohMlpf3KTt/DASzX1hEv3Rd0g9bT3dG
k8XTIQMk7ISNy4sRAl09CYThW/jhNT1KMSUG8ck58jkAWryz10xdMLL1c8IeWMK0/t8XpxdvK+M9
4H0yxmRNHylccW575lWWWBm/5hF8kEJQc4FNRS0p0MQwTOFhas+6S4hb0E8pEBQZXJhYpawmCc/a
0rbfM8ld7///X29+g6IXZ5V6LCUwgYIQqBHHQ/RJwaa/Osoeq1HtO6DFlc5gJ3gB+Qj3OvCs2njN
dNd+ULABqFmlFmDSppTgtEsw3CIebER/s7/10gQNkyjbZlueaGZZRr/Ba4NPd4X1ZSf/KHbXJd/W
ayfXKnD443kaY2H4ikM+h42flUQ7X7XVVwB0iRaR0MawBLentElYd4Jh42WvAQ2qhkxvngSm4hjF
Tl2R3OLnB1dEqvuDLz+yQO1XjqewrkzyeYUcMRr6vYfvgzor8JfQKi2FosvTkhgzv+i0lW69ZiaB
21YokLGbeldCaIB2ov/miBU+qs+UcWsMGM8rk2tWNSXWPd0uQY/DHiDgrJRPxNgk2G20Flc99f+y
Rcvw1GAxM4WpnAv30RUc0Jc7LGhMbF/1sg3rOh9tDj7m3KXO9SoisRU2v9NxCpHVN/PPHshf/rYk
b3tJ2DTLMNAnXXBu5OtRNpaJNp9oIee/aO9Gynxh1x92qgTeWOYv7XX+/NXbcybDDFOmzOcXvYFC
acBcPpk/UpBSBCMHsV+f2zsIrWj15NgZScUtfSaDtcWg/stId0XjYXH0UR+alo+a57vn7z/jFc9L
FOB8UQf/daUORHNvblgSz4i/gpVF6XqFYDiAKg2ymaHh7Z7mro3a4JILDeBjUuE0D8EEekx7GBV4
2ycSALzkZNCs9xhfCLDkdOGb61g3kmCHMOgY72OxyKwQPI/S8Xsteb/vvZAKdgpIv5Rr+qrDdLp4
VfUiTC58Y28oogPMaziLHgAlVFFCfZSq3dRCD9hZW9MzZH7NI8GwH7hUq57tzEK777DDlCyMpc7Y
pzGWt0ufLQtlePCyulzZl0o6XpLPrlJm19o7B9iBIJt6gOc7UUOdQZf/n2MHGYQMe9owep9Pcwyg
97KQnQE9YvLK5Mgr1v/lNGeq9DENV+f9uYtrLYfu4UiWHypuIMlk7P5Nd2VQ3ERAktlna63XwN0C
SpJT5Yist9z1gT2bk4kaVr8qGrhiqrloqwnVMSsKegAwmqa8OKibTsg8C6QuFwtDglkXdeulXmLR
2dJdlshBgUfUdPqYF88Ld2i7NuTLiGdAiGieIDe0/EftR8xlaih2FtLGeoO2OZswq/L3WrrOouHv
h76vpjHOlkT1Wg1IpyhkxnmgQw7EFKnUEQGlDA8peqcn79v8GbxrJ0kf/xb31z5UdrYLYBftghpG
uOu1u5rP+PB4W5ZkAyO4iEIdXQo9Ji3axXFlMtUDi3vd9tctyqy+hM4ruqt9yI6mLUF2LrXEW0pA
hggR3E8zadYfFoJjfxOUG9h0Ex+22Acl65xd3u8oV8hAYrAXTtRFg5e//0lo03kg8E8ZC+uZCt9O
NOVBtWrzg9YdkXi8dGLfWLrTlUpQkkmsRY5/y+S/+ZIE/Kictz5Lk3LjNqEc8wgiA7bhgEJQUbHO
YmjGsPcgJL9COE+C+QS2FelCTNYvjdCork3FVZJVnOmo1Mh90P0I6P1XqwPYW24CSiQIsmwWwrq/
nqNtZUOriFbjwzyhZlKp7WLWQy2E8x3kY+5lXnWtQ19q9sAVW+EBuSLfMzyBwumIEXggAqwVdjSn
uctnpOC2LrdQO4qHR0QRphC7gIDoYRgOvPhq4M7Xvh8z2orR4CaUxVSXOtlr/nV5BhqyTYgacuB9
Qj7nSAyadGp2R/+xDwMfK6EabMzR2uNniBaTKWEKycFRMV2NWXBxQH0Yerxd8CK6PbRhSUGOj4jU
DROSr1oNxoBX5SAbv65Sof6xbCK1mH57fZfYIAHJ337uNzMgtnsBHR0APHhVliJsol8afsTAf/hm
FlMmVK9kehUrfnAdr7L6CP32o2fXPToLo+0bK/0ywHeUN4frJO3ghkCHaARhokoJ2XgDVwOdujby
9dbPOH+s4LQa3BK1mo566wZBBKC0JxS+9CM+/auPgoRZEaA7XxQaw3emCUUSSPRVo5aoXHL+C3Mu
5FepkBjAF8tEGFk3BnVJ8OBeEe/Y6/Uw2+iZBNfj+qVl9BDq8pL++MJA1NQ4O9Blr75UX2DpDwnX
WwNgOEuhbd7pMZyPW5TzSygpZ0Urb/YSxfdEk4WPHyIaeIcR8kXs5x7Tes8nTuCrCpJxEWstCCsR
WsR75qosMX+DU4LSJaX09XDEAaRPaZ2AfJk/7+KXd+qysEiCbqwpLQLCg5+zAC/PxG/z5YTppvfP
lBPRMz4L5t6iE9UPsiQ77ijN7B9othp1YvnnvfXEvU8pxh3fkXgWWfgEfFYKeRkK1DPa0ymw+XzW
OWzZ26pVY7UBACTRiIQSdvMsB0xq7+vZX/ez3ZfQ1ZE+9alOneOVJhczkNv9ba0ro2zTEvLiaFqj
lKf7fp+eOPKIbs75pLGYrpMSKLXr8koxOdc7jl+ErheXKPPwZDTXLLqY3qWOIBJHT0O6v3DRkcCl
P8IMlXCNNELsSS5TQbKPHQllc4QEMfTXrLwkfTZa07klXye1gPf+k4RsnazM+Cf4ci2DhDqw54e+
ccWiDSbr2/rdOVVYSRtOqWRqWB3GkFdePPI7McA/Ol/09RL1T5XKOPcXLoZibtNqtR0gs/fRSbR6
xBvONzBwUDPY2R0Wp0rqlq8fvEjSIbqMiWQ4mnnFxehzqlG/k1dX5KuX8Xh2tphRfKNPZ1+/jrAe
qjeDb0vtZBfAScR4sY/uXhu36ihLirNDrcLoo8FtAh2P9PTW8XCGoQBdwWRNtMSIre4udgU1JKiO
1P2yJ7CqAHp5yvfTAUHqNUsIzBC7eluaCkDlRN/IKt71FiYQfpcDQkkjSzFNI/M6nrNgLRizTl2n
Y0/ZOTo8FOvA/VSTf3z8jhDdlJ4eehTYUAb3MHR9m2CTW6ymyqacLCo1ae5CJi4IkSkJpFKsuLP4
c6ghbCvt1VjUQK022GyLzEAjfoymNdtEETZasOTOlRc10FupjDfDkWX/ABo+peuhnYRbDW7iNqqS
jGKJuVjXGI2nWsY2aVRwJ4GecEvISbdwpFsSs+zUXOvdUd8LRfWxyWmjnJotsJ8f61pqmUEs7ura
iFBq/ShcsLtdyib2r/CATQfR2nNEtF9zaJYn5QHDGAqCFebttvCvewWrRy1XhnQIFPexQaZRBDrR
ryxtFKRnGbzaXJi6gUGJmxu4xeegYj1mtB0HQqEczGOp3a0tWpfVGcLMAm6/0k2h5/f5NVfA6BgR
x2UKcgAkE2CajE7858pc10/kWwL3QQdj7KLRczGh6cblBtfKNmGAn//fWjVybn/7VTnA2A/yNTfv
8MVsjxhQm6T8+YUn8Qg71DpO/y8vfGnieLXzpBW4wjXPmJPLnbA6DMWlJiI/HN0CCvyxIUQLCz5G
fQEMf7Gw4GF9ENGfaWz1g0g8JxjjAm3A0/cV2n23ZrthlMvDUacTo8XkZHOvu3153+5tz2sV7hpH
Vc2vpkESsT6EclLXOBksMELOPbV5MqxLh8f2UipESF7mx09HZNp+2IgXd+10iPdxk+f6XfELHegz
qbRptwE1ejj1wSd8UAGK/R3qEBfGJa2vwTicSoc8fMCsxsW9A0YcHxJfQgqMXF+7AWpHdOwGjS+b
V0i2xbvifwdsmQTWIkRKeIEMz8lqX5LX1vSKq8SLIRlkYTunUJIPocjrwg+Xq0W1gj7msaHOvilk
ISWlP3Z7taGfgs1UWV1oaYajknoDiVTOdzYSUdXBtGBikfAf0kAVcof4DzyYVncmnrhInjL29Mfj
NGSdpdHdpcwvfbM5z7iaEeWqieE7ljys2vMg5Cz1qEB4/6v88DdkTzKfhGB2NTowG/4lBQKUkE+8
ibS+4sT9b6OkOxXzKHrA2j3hZlubV7bL+7PmDs8syfmJuB9QiColhOAj87/FN0aWZahyl+lkHkjF
NNV1g1qEF3p4m2Fk9+Vl6gBdOCxtOSTJh+IQKXBkenURYCjyEdaFjdmMyxFu/jILPnB4dyfVN9Me
zK+PySMvMrYqSbcfZB6uowCxx7SZ/B/8ufIX1EYmnPtOrUCunrFpO9d5LQvtDj8ORymfgknPOYFF
9DqFAlsUFXUxXt3NtdJfcebjJrjxevSbm92VBJWubwJCtn/eE6j1VfRtourm4nN0EkjpVrOmpXB2
HhmtFH/damJQ5dJEzqnTWkLSQHg3DeXCVgWV2MX2uPSS0CxB1UV3UnNi/i5gpSWsRsDKDXMUT/GC
wIzIStXd1D1ac996fcCSCV18c/HZSs/WZQVG0i/kHBlqhqf6fIhp4IPxyxIKarWPPu4oeKpQIBn0
S4t1W4XHbVfKWVas6kAkdFje6F+BWbvDf4lUDl3r5uduO7PwOTIBQWYa+sH24bOPsuCp6n1X3OIg
re4Qo/CXiBMkP7jglX4pnno6Cp1G70v05Qo1HrnRTXXXZi6r1GJI2b0niOhHPpg5UaeAkbL+IzsA
4oNLAh6v/4tKqtI0UQYvn7iSf1w/waKpGJYWhXziDU0NYpv4DAIi3XwoSMxDKAkULr5qD+/Z7qgR
M+wJ5d5hUIo2UbRwb67sedBrr0DSM0J/1tVI5qEErpc3tNS9Bw/4TmORTRM9nU/KSVxhED8pyOHO
5QMccxt+fl5k8zU++D+oMmK4zN45O7ZRbizEH/64vOsdqU7lTDKBGz067GX64DAZomf320NJ3mnM
tBXPTaqL8bMV+PGmsKMDKagklw1DLIgA+4PnjhfyCeqssBRtMyr3DkGVX8yTCllSsngj8R95nIsm
l+tjB/+Pq7OuNcjL0cSEb0TUw4/vgwR4AGsC1OKENODa5BP1+U40CLaFN/1J2WZvYsjiw1zJBUX0
FBTzSTUHJ9zxCCkD+I50JS0h699wFkup3IHuYO8/832gE7J3BvqGU7NVArxlOljKvVF3WFvXTNiz
UxhMJ+fd9GFGc1Ef4GbQucud1zS+rWRHMpaarJLL7z0jK+E6TN+G0gKAWX6oGeaq/1lBBNWFgrNc
VzygpkzbXZ8yU3sy5fzlASi7GSYiODk87eIXtaqYRXZzWQPhAGL3JXYi1R2/PsfmjJUfViL5dnu5
unH6D6NDFg0h7AcABSX0xdgcdxR7JlyiPBMJ/BAtOEck5G5jJDwuoMmW/MQaKUE++rOEDm1G+2dp
GIPHOZXuwlOusdfKMiJRrC0zIbBhEz5ACfQ2xtkUZeQuVjUN+7RCN+ilD8NZyVmknnAUqFS+yc1M
cAeCji6ZO7x2YgbUI9ItZsFB1WeohPgRH1cI9k+eUYSZLgoCIB47KAIs1C0pT6Bide1n+ktrKu1W
HaCqANNrWkXAy5bYSzCdGa3242ZBftkrzycFVYihQChxCpt+ti7C7tYRPye6d9H8o6YRzie4Fwso
WGInN1cdGCAPoHQ5G0nVxoIRHj0baKy6c7pa9WhIhsu3rYNzGzseC+5Qv3PF9R8todS89AgYs/1R
7Ba/sLyWqBGYsMUcgyk88DjMfFtfCiPLA3G3SDBvEQ60DjEYGocmKCgJtNokVGuGiioR1kI/ndwB
B2urGzUUlDRtHj3u6DjZQ8fuX9mGq8UcO8uokmWgHo6ms1DxsHMD0DvNRA/OquHt09ui7YAbcqMK
MZ2+tEQgKS9QN/VYuYjuQbdbx+FLT0FIWiFKDK8TA8aId+pJANAuh6SgZtq7VIDpZp3WyLqfHP0X
ABFGmMur9U5TMKqz371UdmDy5AtR//CaC3K4q2C3Qu4nTnmRZ3XzoL25Tv1/5PZFQuTB6dppO3dL
oeI6vOm6hnoW6hjR4RVITfHn3wuIA8Ek0am3nw3snalLkaKUNp65GtTw2tE0Jvl4/9fiCL1jZ8ah
f7Pjf9zHA7jXvdgWLnhkl8yfJQLjpDEtsB7i9b7BzQCHacQmzb6dBIawzygOyr6axav7IWXviWP8
kfX3dyvOE/vsjhK7rtte7yiFs7YGORdMp1XCIQxeyHDA7X4tlXbILBVInvYdIJ+2YgiOYPIfLzyJ
JnajwxJl956KNcRY+1HplOeMLllkk+IknMOuUXKDKDwODDaDzNPb7X6+7hYmm1kjBD56X0E70z0/
jO4c7sT9yfhjNNTBubAMZ7g4uZImXKyhhGpioBZXmywuwqzM183av663V1IYmFY6KsFSGU5Q+A2B
nLwph5gMMdULeLqw7kj/j7JtwEuun/vfsrEUgHXMmsdHK0s7zYOd5PZyuIJtEsVbkklKhnr4ZqXe
yxZcwWiYBxFabKXzyjVoQ1TwcoRZgr4vxSUbricIic/H2vVHpDZYeOTBp2xjeUyBDcLLEYiT7wzj
G5Vg1APKD1a6h7MbghITrioBmzi55MHGaWffT/ZxvXrFrdsDlayOLjcG0PKtreOZm81xUYWp2V5Y
8Ap0waAXAKypQXtb7kVshKfTN5k51N3wrtMbPh9kb2VY+nqFSvewa4LzkfanBhN/VI7IpzCas2jh
/UH2opiQfdHAjdRBEBjoaMLERAtxyEwqqc7iHVRPp6fo+7hm2VjFCCV5gLIg7o+VGMFw0dyfixDS
mIyj7CUHJNpewZsSZZzLxDQi68MnDaKV4szoaroF3EbHIIyZE4O787ih1gIvhU/t7kuLOkgDfntf
HYnlJ9YiFMgHNG43xDgViPA0khbDjf50G9W95h4xY1rAxjuhve1oewgmDyS6pNq8It2B3iD7VSr1
rDl3dXT/xuWCIFguB90kfIL483v8KrtqH7qryCN5g0ZLVPm2cqM2yCsuy03wxCKSh/kWPJ/COxiK
LY6Z7xhGz11CzpOXcOIn57xsmRJg4TSJ4PzDQeVIp35151vw9I50PkuGEfoLCjIQ6jl1zP7czCT2
LPGrJe6sAApzDNDJU2uqV7wV8I8EZiLUvR89Wd+EpKfq6jmmgwaQtwx6mtS3/Rq1TvfLEQfWgZLQ
CK8EEGZb2doDh1TKwUyoJelnxr41GWig6TptWczd+nCNwq+FZZ9NgXo315sWljFe0X5ic/hiRia6
jnOJVfD3penrc8eS+cMnr7g4w5pHHnYysvIGAGB9Vc+cAY6n8heI3D1JfNj1GdDJAe1ANn5pePGx
s3+A4DBjBJi0XSbSWgFM/10OXBCHYhfkBUX31nxSDMlj9d3ktcqqbGFwLdoJ9FghcIco3KR+sRr7
/2iGINpoLwO6cA1b2MzKiEAsg+yedFvYgoMOC1Upmw6o5LhqMBpcdDmILbrBLC3X5tC+Ba3u20us
cU5YEgbvsHbJaIN9iA/R7XGI7qbtQwVIpu40i6RLifAYh4bBqZfMI6k51Jc45WkiYpj7vIq6DZQj
HSQQ8bC5jVBOYGAB4ns7waUJYOBvtTpl3p/ccJqdCosKPCrQAntcQXRi7WICHOG85aruDF9RjZW+
aAat9dH8Vn9qFcovCCYKA39vPqjwbpDeZKgw5NlfMQMILrcr24Ronv5jEmMwaUXJ1Kr0VsBrcsvA
NX/vD2H4DQAvDHAjBH97etDlUjAUm/lqdNSVsL50o08A1WeattANomrJAorJiN9Vtr40oGNYTiaP
634iPjRJit9jIspaAVbPu/2oLAEArYvabrrFZ7CDlCCQc7CMY9GV4yTBTj+dq54ymcyarmqh4Lwh
SawFxkC+fN2ero/uzxUsJ9CClDcn6qincmkU0cm5CwFcVgvF9ICsfjnClaoogA/SEcQxqHithZfV
tZ9gcP25ZBp44m1U/5+jHdfsqa1w/P0mpiCqIiOThyJQ18ZoIo8ttIN5SMUCcDzGjNrKn3lVt4vm
3QSrSbqHOhc4u1+jCC5Y6qsxdthSQ3B5hBAMALYIpvDm+95BM2q5OEG4hyjxMo8wqSbWXv+ifLO4
pvL+YcJpvIeLxmy41hS8fiulOjqpOodMGo3mUWt39i/mwffiIh18174Ez9+32Xf1XyLyH3rwt4sD
E3SWvd8TrIQV1vYpeJonRQaSzS3cNAEePV7/Z7jWsn01aEEgMzv/q7jL5rdfaZAzup9yupZkK0y/
ebdlbEsHAtKf5PXh9bxBgRcyrRMZuVQC3qDsjt4JX1hcSajEu6SLdAjYvgNTaC6YTNop59wzyN1K
IG+J8B/t5iyTRyHj+M+pf6ChQvRLjKrrY+E+QxErmyDLEzjpMO0iSqOCNAcj6vLKQxikdHdip3Dp
vj70a9cPGV6PFlgKMW60oMY5FfvFqqWGThmY6T5VuOUWqm0WeEUEgXUg4p15SdOBKYH8jSmTrlVb
P8wOFoGZ1nel1utTX8LjdfrMnL5ZtN+EgY5f+hAcjYNPMVyb6uu8SNZmnCAtWFC3swVVHMqbLSN/
dg/WG4y1IPvCyuZ82V3HpG6DU59rC/2xUA88jsuhitgj60w0E8egXJ6F55ZfttnIbx75MXpr6AcC
BFadf9WuQOTQZZBdBSKC2SPhRo0spjLGvc0TVktkVbOBATqZp3TxffE3g5vc9Jmd6oaSVK90Lw2W
4dzhLgApLg+4oQ3Kss9xB+oq9hC+EUN+wx4hJ9J2XRGSp7iguCrbbQ/PRSbFWpk4TagVmj8wA6LG
XMZEmWkeqOQVLOGYBmx+g2+uRm1Z5eithauyQ0FRFJP1IdNfWucqgU4VXCGvsvTeApUXkLVqV91R
loQ72fHg9AmOpYLoEC+SGJ1NkVdYuDHJGPnjxNMhuHi2B9l++GSoTAyfnZZkoijuYDFPMy5dC1nP
4yhT2t5XEoJ7XxR9we8VYLpFcz1bPy2yrAmtvNSEUL0PVC928+hm6niYMLSymV1WzgkTH7zNMNig
DvgBTSHjBdZ11xGUKY7810/tX+juriM/6z6amPga/teqLlr+IzvXAZDbJvcItPX3qB+jFZUEsVpG
rXJer+A10K5kMADuslmLlQgHe2otLMpJDNzFZnXNEn9tQL+Ve9zNU0j2EbwLH3LE3xT1g2lknIoO
RQYykO1fDOqAGGpzW/c9l5etd90f4TNLqdYhuPf5kVfaJtu6XKGgJ0GmgZU1xZn0j3aXc/TFzEZT
VPtuyrUMc/keVDwnNM5rEyRT0vxlcUQrcC14eUlK+FPuOK2SDkuP9NqRcx+X3pfVYb7EFX10Xnse
Zasgs5e1Kog1zkZeqkXVT7NTg5nLLeyiSDvUXOJ325NUun2RNRv2vcNxY+h847sw5gVr4gTBkoGE
J9bsWall9hAN5lqlACxIHUIKrbcfT8npylcOV328NWm9oVIR1GlNRBSp5S9AgV2HfCAA8wYUcgAH
UWUnCxZyVcrCgjs1qO4SKYVAeIHrPyFSDB2YcynOJVNIZ8j5VU1WttqwG0eoNtwuv++i8AOdXxgQ
l7n2VZZgVG+vYyPo2iEOVShBABh1+B9R+yngv8OKpmnIx3GhFYyTFef1du6PbPWixxK3+anotg1d
X5skMXq1P6yvzB0U6JvIIQCc5bepXefc+jNlOFIgKJuHq20ceU4w55+ZVVMSecW9brqLvMqyVJ6+
I0C1vS6749bRcKHcvjQzvCHcTZmEkHaheyXSTKdZDIRPKiOIT+tU952qNdguS+/bBNvjad+djudt
QvqpsNIb9Sxf5t2OzIaZItcx6fKjLs5Hn5skT+lICLB30l38qNsXbwRLsRu7CqPmVfwkUyhzQgCU
7fj87xgmN7BqjCQYNKFiyyVhJRsZrWuS7p3kL/0ZvYd63rLn5xoFT0As853uGDF2oTUdptFDcFJO
Y/I86RjTBsXUs9FgIrZ3NnxnjICsDW6bLakRqL7KeZ0eh3mu5wXOp6nzevaNk9nZnXZnKaUnL/Pa
Sk+CJwGaxL09qsYlSKFK0G2Dzb1uMIfPfhh4HxuPAjU1+WNDP5P5Zx6cELsFYxlqOLRPthgYMPtU
UcNhqqk3j9rlWN5aFIs3nyThyRFO8wZPWhXYROwZjf9hiBhwTfj97kN27jv20P4hnj7KyUqBxJIe
cIxd1QnqBKe/ezb1B4wNnjEUuJaaAB7J+a+lNwl04lvnl+964nFES8rkJ4Nz2n5ou+H1PFZZLsWY
KVzYa1Tf5MX2XHmy3/57g/ITIw2wSK2kE9hSfvW0CWYvKvt5kHPxqBNHXYM4CNEaqHtrqdJOHaNo
DeciicGhKT9+8jPsZCbaJ6/KUm1Qtp0Y4YbHbt9fWtvyZz47+j+yibt1sfFVgGCZTE66XtR1JXFz
jTj7x1Y2UewSXoy10M21UShVMbRb5b2r7As6oQ7ZxpwELNyB21kRQyMHLjOIj0N9Mo9Inj2m+8p6
pZfUvf9hYhPVxKN0qlTAe6qZOFCzA+TcFeIKbBaTeITTTB4/HcJSwvRGOBPKya1xNrEbwDcz1ee4
H71r/WkkrxW/gfPYNBdJvPBBGScxr5EX778Jv8n+gubl1OgOH7slV+17VkRdKyIeW7CowGJE9F5W
BfG1nDe/NoPw5X8YVmQ2UvjLJ4oxZ5pR+iYe5LWSUurnvTLz94UnuUijQq6dzYe4vbXviL+MsWWs
L+DZCYWRY/xl3G6NOx3O22fjXlDEzfDraX87bTejZUF/c6VMT+XYid7NrT4IMs6neZbmFfX8M7rX
OSVCSfIjPmjEDDFCAhoB7xV/P8v78nZvja2N6X6igx07/sNwfXxmT4vjuIhMoSj+m13DdjejEZO3
5FUypp1rzx+At2/fSwESbJhpglvfpFp1WrQ9GWbiApLkeml8DxfzhVjv1Lel2PG9uhL6FxgGn9Sm
mVrzZpA5wAgccktW5yvVWKpy/Wo44uX6fAHjJElGsG4FnjFtlqbbLDJW+KONWGATUJ11sfgrQAdo
OWc8K3b/7MLKGCjVhM8C/rk/vepwx7ZAgmSUZB+0ufQ4njSkbk6UXEmV1q15zGMw38jghgEdOw8U
lDVJY92joQDIXzg/gNnHX7APP3vwm+LpinUmKlAo6SOmA5EmwyZy93Of3VTpgVncTr5vhj0NcPUl
mTxwOWFmy7AxRK/ilcDa9V4kNIeeFZy8RdIele0cR91X+FFRI4bzE/X/rt7IGWgNUPb/Z5Sl4LIo
6H1XbTUF3orfycoJTqPWoqAmBDEeLaN6y9tecOo4JbgzcD7Wd3pcW6uwpl7PAFWdPbrUxf0aJvjE
ucySnoNwtKiCMEVBpfdx+zjR44yAFFrq4tbph3YquWiPW9jjH2VYDSMjcLYgbBACdbboumw4Tlop
O413PEXs29gID4bUqL3x98zpBJvQ7t1mLWLs9Xbq6lvIgkJuPDv6gUw7KgfuPaLLfdSpQvTbuVgZ
5/Ih91rlVi7Bp0xkLC+SxfereF5VHJzuf5P2lLzz88hJcPLMD2DSC95LveFJOCK5Z8Xb4mHAdufm
syIu7YJWLw0qd4H87MfW7hTe0huq2aalHx6ZVExuJ6KwSha/SCTwg0riKMkY6FcT5kkRuWT//3Hn
5e39URz3tGAlVOvMP6VcRIH1S6cde5suziJuejwP9MIcDsvjHS8mIa+Hnvc2aucbWBqsUUvCZD/0
ZF3A7XXx46386bEPogyDUopvtSnM1wCjw6k5v4uSUUPqb8TIAuRK8dhRal60NIQT6G1XcsZtU/+z
NxC2qWBGwlLENqzjq6kiWRrdIWcr+WJ7b5tP2Sx+T40ElGvJDsFeMH+MtJ3jchHgAlHpfy/ns5K2
kOpLR0DdM0VXLUdNhZ1vLPlsTAUmmD/z6d2ovmIKCH72McZVKn0v7fenQDfQBoFVS4aoRVBdVWZH
qC8ifhMzz7RrJ2ciT7OsV3mqvyWg+5rm8DVgUds1IsbHMtSjGMw5ljTPcgQGseuCXhbqhm7qZkJY
y1JmIm+n677NhXwFMWDQ84iOWVP87fofdaWfgelEasddbTMRd/zl/4Ltyeg4O4dDYnHN82IKCMru
DQkpM7Z1OhxZPycKDrsNm8VpvD2Rzll4TCxEAiNdUsVP0wpccbfOBL3Q3RfqHj72xa0B9qW794k1
wirKwQ7GYLQbhboVsw3aSpX1y3KFFdwljn1P6IBdR1jIbw+pS0TeByHkKXCKTu61yhLMljazifnf
5YcZGjwwtYKaDdwmDv2/GiimGEeCJ1fhJ9z3oSM35LTBuoaR1JreYVpNgIlL+x3+toM3z/bbJAe/
KGKZb/ip9gOHls3TmRvsbQbgycv0wUd2Wh9RcljudVp3zKE0iASjFYXZS6hifmUpQsVyruTl4Bos
ngthBI4sOQXLXdaxLl8rzIyNqH3dl/2uJEYEsdQz8WhjBsUEhEYA3fFvPmsrAh67Xa+wgCvHRo3W
zEMrAERPBs/cOaH1BSMdpkbfbaC9NLn6sBOzYfVTiziiucQ2vWPiLAU9SIrU/WpRi9MCtshNy3Dp
IPTNluJSh13/8Wt8gthkKswNBBZ+CCmn8M2y3NOHqq09vodSyGPrj3W7dJF2eCs3c5dyvByjmuPD
Mn0imw7Kk87sMuafPtbIRQURQXvP2VLjTdCcRPQbevBIbQ7QRhx9x2da6KDeXW+ACugZmJjuKE71
TWH/qW6KOkEUg4aHM82hprZ/fH0cfSYdo5pHFlBwb33IxZ9EwwX6nmoJQ6JCAf9ae0g8bs5RPweq
SHSKaNWaJWW6pG7wYPuHsks7Px6HfXeEP9daQBG9uWAr9/pkCjd9v2KCxwYVmJnt7SLPOaCn00KZ
G/VYAGcoPtvIAoaSp8nTbAVrKF0vxkTGGwkXL0+lGgquD4XzZmvdnZVym5P8qqM3J11MYXIECktM
m9uBc6KFZ2t2YDwYQ3LCJf4eHXorxNy6mjAfkhIZU1fVgyQDAEnJGkJFV7dApUTgn5/ayoQ0CnA3
4kbeoeaHI2AxIcFMm2jS8iAanNv2jLIWUdzWk3DovmsK72H4eo/FN1+5c+9RhE3J5OTnf63t+OOL
YnMWoYVigzWLikMbPzkkeLZJ3DmaBJ5wiz2lKtfep0WfWctu5+hH8SwQ5pzRd+PTJ01HljKvzxy4
m4LgNZBHzdl0Ka+H4WH1axF2eU0vegkSgNrHQpaSrL9zCcM1xvChbkeF8Rvh+IlBW1kTTvgaop9C
3sML9zyy/SFXYCh6X6rI4q/GXQyNhxJOxHXRFzxt1ecocL1gR9uc8ddt45E447FwEJGAkxI3FGaf
IDJN0wfpoCOoOfxRgnqGqWH9v0t3hEWH/w2GsXdyXeF7Aseew0cQQnbKANwsBEKB6d+8EaX0Ytnv
2PNu/dno3Si/VDigBoXYrdF1EPVnGsyTGpRIijT1cpZY8buLw6j175amedZx3IjRnmZEJVL0W6fU
o2LK71CADO28MnwM/HRyPZDX7Yx+NlkC2b8rxiPAs0MhL8upiO3pGtOoIv2Ubl9KPu2RAyRkyxxu
0tgDCU+gnP03XDPCTO+F1zTOSMAA71iXyJlZU5Qt+3uF4c8Mz1BiaU+NEtouxYUyy3wvh1x+21g1
3/wIGKNjdbWhIYhTxC+cbwAKaBZdcSrfKJM4VfnyIRcUcQIWglTTZjUsfFWq0gxhjya2JbP1KZdl
ileDyTGuSSe55JhnD6TmJREoSrCWG/O2W8nEMz/81jY3tf9ACACxk9xDfmpfDUbf2vEjpiYIinq1
a034J1ssPJd3svg9NGbkwcyw11P8QQTPy40ogINoVkdjzFR1pChNwd13QDlUfqPJnko6UyZeu/ML
3xs51JDYyfmPuEPN4Usdv9uwvsMfVOG1YTwazreD0kksNsFHU8rWzrlglmG8EAQsxScCEN2NO1ZF
zU+pO3ftAe+50/K/HQu4fMasl4iMKULi/POWcL36BuDVRTmX/cY9pZPfekJ1w0YSYqYjK2guOoaS
FLpzF1A2wQrTAedGI8oGiKbMKTLWA1kve8TPDW1O8xCr9BXMnzLl/DdUrD4mbi4DMwQ6AfEoOV4b
scyvCNobZS16965ASOFw4CsdJNAlLCnaktCbGdzJmL4XtWv+arxP7MXOndCDGA6s65mIJX3iJh1r
l9ed3/LwF6chUoH3gKcbJIGHxkxrjYkYncQSrVWtamzOCsbdQ/3ImyjNIRiL7Ka+Jn/gkxXpmWt/
Oi2WtYjLBDgVWOatZykSUUSPwasG4ITgm5+UXdQTOoxUvEOMEnhHry0webxB27Z8JkOYV6c46In6
86pZ8NoJc3rNy0jqZzStYDkKqhT0hf/KqJwgLF6J/Yde/dmWY8j7TMt0mMtwo5+okiVU3AOFmLhy
L5ZB2JjEcvDSxjH6r6Wu2PVNkH+W2L1E+RslelVVNhUnfSsaW+2DouCY8FL+6zKuUU0/srQQPOCl
RwjUIc0qU5jEToTe0v2p4GvOG0HZSuWWnBzz5H5o/JXMQ23MN/rILXJNcDpaqNQu0GxJCjxsED+M
0PB4xpXRKDDhjTley7gp+cWRulrMARUnuofMXGzGtCg4/gxgqdKUH0+8/GJGyWNvQGH5OOeZrYn/
fHFvTboW+V5V+Qq4iZOyOCXB+4EWjgp8L9PcRxSQE/pV+EFRJBoavami3+xi0ax9Utrk2TN8gQ00
YQEerjfbF+Esh00nweYxf22lAaEjwT0RTRgdy00Zu2o8Izmqtppf1hS7Xm6heLX1TYbGiG3CZ0FA
iIncfjI0K9nYaqwj7dwDE0JQGI2vTCx+7kpo9GQqnX0bODDBsCeh6vqTePrQinb3i3Ll+00C0x9z
S1Dyi0AB1ZVjkjpXjJRmypSfvykyKp17ELV7OB9cM7L7V9Vl+vczFsWQ1INfCYsn0rNSPW/zSvUw
DatqVJXzeV39baa4L5PTrvFefy14cfLrrq5Bofe80FY3WRb6UpIgTsTZskWuYmIkT5YjDelcWrEn
qEXHu24AJyci/bxLhYgh2SsJTcpR31x/enLDZ05bSajuLlHFF7iGk3YdLNHhXOM57IhyAmDKuPyx
hEaGLeCObttxdirX/7BcVSi8Ie9SEo43W1vDxFtgMlH7vIeTwtStKW0R45l2UJm0A3ZveDrPPLSE
fesQ/s2cloPK3Y+4K6aV5N7Qj4bAvLQRn1IRpdH+/Jb07Mx/PpLQHvYBpDXq2qqCkZZzZub90eRg
xHb9wfruO1VqFBG+Ux6ibJXkag5x/TgMI8jTqJL8BAKnYF0PaMTiNS7/BqTY/XvFrJn/t+0xPB3B
0nQenQkHUE2DaBURfpTnzz13nDazwA2/y3BcGRWBIGBpaATEjwB1frkUSBPuPwBwMnU2gdCBQauR
i27nyqDgfDHdugYeQ5I6Q5S9POXuO3cO5IppbD2Vctz9kr+uPY7sIqgxSPfC5TYEivpH1CX07k31
eTZrS0OSZ4JfkRxQMfdSquCRxC46QGZKh3yIwz50pBq+lrgGCl5nQ91fk6H3ik7k9UMkRhttdUJ5
oAS+vzDbm7AZnSpq1iB2zcPSVPxIOJgo0YP4s1qdaHXCCerQLGPRfYosB0aCMrHP9nHK1SWkGpkS
+5yMDB2mwibRZAbRwVrJ4y1Xf5rbB5AitrwNJFI/fYJ0WfLzZauK39dE5id2tCRMKbAASEkIPSKb
2J44B1ZRxTglVtsIQwX8ehbQ+qabUUR0NUl+hawgcrxc0BlodvAEkarvWtglAhE3Fnswjvv1/Wlt
6R/kZ+QA+uS8fbz2JpMl2+GwvF0Ca7RyGULjMmOwkLn2tSEf6eViAM97Xc55vnX8Hx/H5tysRinn
4JTXAGy6EVr+0q4915crluQnLHBhhfa0w/JM12RsdNecLg0OpE05FjP616TV7E4DWMgzzkY0kFMF
atonNHWSoILa8JYKHcUP3lAT6FWi2YqsHDEn08pJN4uQDfwI50DiS0+jWgWTnT7DLzUF4qPZY7aA
iNv6ZlYyDOl1FNdtkUw7o5CXmmpmTvzXAreZ4evgxdOlF1JhXnBFeU78M01ZZdNT+D9b1SKKy30l
l2CkqsTB8ua3rytLkvUCCEt9hH9Axhi3UPma8VI6uaadk+p44TyhQhu6OjfguPAbNXBmhynlJiW+
hqcSXThEPutx3c0DYyN8ikFoPeNJQces3kClTarOD01Pz2XZd0y0fdJTVlGnysKdpiDGQ7ceKW0p
zQjdJbk0CObgpCLcfUnXxuSs0BH5FHlmD5bVQW9wXbndiJyMMQ6gTp5Wd6CZLvU8Yr8HjvLOxMBK
OHnMJzk8nx1awduK1nCDEVVU6T0YmBXwTw0bJO84wYO+pQbVtTGBcVxIAP4L1QLCG+nhft6lvfrS
mYgjzqGxY9Tn73K3cPIC2HgqCulL74YQmonOlRJAytkJywS59dfqPUXqt6VnIbUGt71NwdSYOARu
dm2fYbRXmUHuw89ITELnR2lsxI5K7MRCrA2NFxsCEIhyV1labIjcyAGMm5l8nrGR5WmpqZ7vIgsX
VXNB7c4GwqXfJlpKR0MVa7uaRwH40qUkPpss+lPr7fkCd/y6XZyi3EPGWyIjWRBaxf/V+D1Gwqi2
i7x4bNhKVddcf6ZrrsPOM97KQmSwunjCoV0RNrjMx9NedKo64p0N+QiCflv1B1aPveI6GIveA6k5
VQsORL7ms6wuywPmV9X+UPJRKDyq6GOGpm6z6vUjknydn+UawUki0mDyU7ryVLUv2ASVnlZzCHMA
c7jk2RCDg9fpuzivpoE0ORZbANaO9UgiuJkchqukHebd7DnBy6Cm4xeEvkwUxsdUpPGtYRgUaCO0
p0s9iG8nH5xNF/O+JpiQ+7AAjUmhs9mRD8qCjLv/fTTtpv5rWn3x1aWhCraHuLbI0Ahf2lEYqnM8
AhyIVVPPi4riwpxV+38lz0SFpQ57FspT5DSvfb+V1wfaeAveGkK+nMQzN/jotfG9UTmpHl6Q82ry
J7j2bwy6kP8iU7wpe+WN9xRFRzOs2i2uc4K4EsMnihsnzv/nNM5RdiyWJtvo96fM38iRjFS/MQCi
jRVU4gD/6Defo+OGMGxSCBpYep7GLFhRR5viw3ifgcPqShizu2BqpuH2/xUvxv851AuIfMFH/ejr
K8N4noAsbR5I9t01VMAviQ8Bh549n76J357xByBN3S20mYSzDqnCl6zi6513vzBFcDWuOIbGIx0b
maE6nRxdUSfttmzckxENoCT7T5oLzpErqKcOc3iIihrLe8BnE23oKtA0eNQ/QedIjOuApv32YpjS
sQMw33GVmdzwPenyRIuiZz2up/dyYxKGIgBkZxnEIS/VcajojqBHuSjYHpSzqW0Xxi5oSQMwU3VQ
BlYLojHCvx0mc92pb0popwJK60NOg3aoqUreiOuYIX1663WxAzcVQ2QA6+Eu8ZT+o2ATjL1hN9yF
Ay1Sm/0bUQxqkGof/DYbGxsYtZ8QLEONJPwg3iIFADuxPhbuv+jJt6x4wm3k9Xqvm6A89zQe4gpg
b74qxH6qa5kdNSe8h7ipUQJcV1yQ+pAFjRduAnCqaSIlU/RiA6cDJc73GJa5VX2m47Jyi6G3dCMV
QqBaKYOR2CVvdNpScqMKesZA/d3BrZSE0v2VZSY7WK+mLYCNcKASYHnCATg/xC1k1zbbHj45nWyB
p65h1tDtBUcEQ6s1CEbtKZ0wAW4+C4TCHG+GAi/atiE5FKNWWbylSMXoVQD3Qp++aJA2BwUJrOIO
KoJRLB0e4Sel0GaGsBtyMI+vaLwTG5tO6VlVOGxRm7Ira0Qgf251LVMZCVIHd978M1HLQp+BJJ3x
1z+5XzdsVe21vcnYYdVICfYf3my4Kd9hNdkXolbidSKGMDblcD45eJqQKltTFd6lstdrFQwKX9nb
sCA7z76NLXINWw2dRlFwWHdTU6uZ0Ty8xnlsZeeqYp0dDGSZygDqkK5ZusNTB6KpaCgcVV9wHu0Y
6qt8JRyfYoMRQAtihic6PNuXuf5IGbd755KXOoVgMA0RQr+cXftVh0YlH/f/+Zr+0gkOfRTso+Dl
454cNR6SKq+sQSZdb5o1YL1+0HkJHSv/BOyHHueMIHcn+a3wMefj8qRyaOS4sqgWcfglej28rSkU
eg5fqqMAKcU6x0CHT6o/6a380Rb/lIaX3eTCwPgc6jWJEzMS5yu7Q7HJwKi+LBJ2260PpE7DZsW+
Cl1Fmz0dr8qlaoKgeYtr7JOeqsM6QDUwYSYVSNsT14lOzT2Z3YRNl57aZ2luiaUr1agLHBa+5ZNx
5y17U165Bn9t6K4A/x8n/Ni/so9c99Q+moKv2H+F2kop2YI96Bax9IxVS+T0N5lBqZ+19oH1fdnc
9kgkGJ7qS05HGvEAnpm95JxgxAG89bpF2Ou8Sa85utPY1W7szjW7q11/FmgensUUhu7fhDA4/0Tx
Ve5gU5JEfWSc7hUbso598voiavuUnZoa9OZ/IcgFV/kK0Lfxv+AfXU0GAGMSfnTq3bms8wBZL0U3
big1BqZpbHMpnHaS1I4apmYc69iUZnVlJ0L2S1Prf83dErh912CF9RWYEOAK5BjOnS5yd35vNv4/
bRmow+jh1Sp2KS9Xq0EZgexdvwTj1uHIASeULdUdJ7aMoMt+qzzaqgLjuMymLorgxuAazHPmv6+z
YrNQxuv3SYy5e8noBAs5gWpPPzlzo34SBB7oteeBTcxRhZvii+mAI9uGzjJXw9xwJIwD0A3tPsLP
klCDIzM3sQzjilXlA1GFjEpcfULtRJYGwe03ddwIZmqh9CwrAQYqYF+HVOYKDmqMKyDd16ZzVZ0K
WibQvT7vblBfoF5t/NAIZFAKDpAuqDomIeWCp4vf4e6IDvGAcigE2KD37+wMEQmqUQ9r7LSacUvE
3/+b0y0zAqj5vCeFbTqMM7ywTYaFCYxwY2SD8rhMDsnoxLyN0ZuMXs3biJNyGR9LdSd6fCYu1J5y
vyHMjbGEYd/A1lrSd938Wa7gnPyh8E91DOwH1Q/LKCionN0IxTWwrYyFdflrgiX2wsQHsVYjGJg2
u9/VC0kCziwpadjzSBKt3z2uvZu0eNuJp+YTXBu8mTcWMrtvNZJHTQOPDbiMooEFUEFga0twML/Q
MjREP311s/EG8cNfwUHkq1mNSMnB6nOimYmcLlawIAz5hAND1CGoiZU3MRmc5FZDOw7p52RJetEX
qdnSifBy3PahprjoKx5Lzm4ixrglL2VNV0XE41plfbxrBPOo1y9Xsw+TgH3EbjE4iLIwUtZ/Kj9a
2wLCk8ZktK8o3ygECsbpkGMysGelzj251FcgLtKJIDZrgumI8l0owGkatchxmQ86hkcUt1K59YED
pxEAaieMOMC/P6j/FnU8wb8wQef/iYxJ6pLSb+ZGUH+fKGEChAf4IFgRwAoPM/sMRIQHV/e+dpWy
EHzzRRvvY39lPgpJZ6QThErCitoM3XmLHh6rrdVIRnIcrtCRTCCiZB7y9vzJ7MPlFcXKDxwiO1cP
e9TbqVQYcVv+nH0MPH1ATcEJDxmQbFBmGyjF8t+UIytgbEx6rOn4S9QrhNPY5ENHgZ1ONizJ8ebR
YZo1wnSTaZlXex6121wX/NBBHwMvFtjbRiYnmGU4RZl75JPlo+RxJARbHS1khj2SJz0IxlzARmYk
tKyh0GiENEJPxe+HeJQWy3ZAZj9r5gLWSvU0QOnSUYwkg54vNHrb9tyKGmGRu6FkEGw5ms8+BZzW
D5HpE1UVmsk1cBWspJkrlqxRP5wd56RVXHBpaINWpkvxbV9zhodN0k4y/Aiu/PqwzR3hTkB1IO1n
pGAiFTYWIPUkBCBtMBXf+szius6scN3xysSJeg2XZhyglS6yuyiqQuoFrwv/aM+wRvyzu6m12VXT
P+0eJMJJC5c/OVQ4aem0/2cjEwIDyQ+Wi0uHWkIxFrvKZWW1B6K+tmY1mC3dy8CB4p7KzOX055ed
SHQ7i/AGUeuRk1TkDnCgq5XXBWKMARDNLEjhlM4ZWCvb/b/GH971pdmT2VdJUM2TFFVaXvs6lGlP
PYyKzq/QtLS3eH8sH+Z/6GbOEExEArViRX2Xsl9om6HWHIDHSLm3S2NcIumxjY2J1GxotUelu8Gu
T6vugiXgxl9CZWMcAtaIJNtgsO7uBQ0AdarWKT915wpCHI7nXlJL9IlB4y1KWrPZVV91LzdXuRAZ
vcEzXodpNed2h55bH8G1WQ6URA8HOVH9ufqT8jLci969ijc1O+Zwn3AkGXwl57Hqc3E4eFDRqhw3
wHc/+PhqHQ2IbOZwlMHVCaSadgMb610ZoaqRevOC35yqyr2WLHzHdmSRGVJciv8JKxFJ0a1vBVmw
NhbMjPW9u0a7gFao5mUIEDUMJAym3NxiHQsJjrMHce4+D3gHblBMz8RGZ0SNUmybknIZsLnJxXqm
9MdlyjRTNOMOO09KcaX7gtMzk9skxE/cvIySKjMv6/PaDSqDWdX0oJtM44NebZYaGd8q9nx/+veZ
SH0OAjsdxIecL/NpOjW8EpgvcOfF1B9EP0XaLa7S+GvJep+8oWJgt0UF+EXfXQX+j1IxTe1gUdUR
VpVAU0a9Svl30F9PHDkCGcHEmeeEmmSu9Wyc8Wa7luYfz0xN5HRoRozTWHacR9nBMXO9gkJLIpsq
0caUejX/r6QSeUFpRLtqAmC2NPq+FBQSzbCU+M/uhdv3udhvJzNWVvmemR9CWeAJ7M1fzdU2z7Ln
gOzJL3OkeiCASzzvm/dk1MMababONlPJSJ1JZo1QM8HGR9TYEATaTxcuVVFRCO8hZ5b+sm56OlVB
yFBR7UvWLsANqyBrnBkbWoxB2C5OoOBevehUKyXc7zf9Yt4tpJkP+fOzqhQZvJj2Z0kOfB0Ng1M2
tOe0+lmabkqOAtak40yPAsayIv892dK58o1gB3ZiZJzBqcW9onyHXuDDHWyETy+j8CJsENqRp9UA
l9lOloO95Iqu8XQZMn+8YtgIhJElYd3w/xL4TC0cLb/djU980+sfhrXJCAoG5FMeSBcO8wQnEwcZ
80cZ7h9+0zdvGQYBRVr12AUPECdYIW+3G93YmiiMHjVlSuE2wOKsh5kXQP3/Ogt5IueKgmwr4tUs
23RWlIBB2ek8h9RFDBgst79POIlge3OAw5R+8jhW0xMxvnlmF4B+dmMgm0Jr6TBcS+LnEzrOxmod
jTik+ETEH/JRNz6sv7Vmx0/0Nyd20Gal7xz0/tfwkwt6ZPRUpKicR7d5Wahy7mPxUWRfxy7386vl
57Xm36DCobpfJwDmfp3MV6dWBDoKWnaRSTFv8QVRJdKvqObODYrYbFbNbYLRHIjewMl+e71acTbW
Pqjqq7eiW+27aczUp9fAW9ko63tQlpGJmkyCLnNzzbCZsNrA87i5NT5sInIDIVvysF0FasvYIsmv
LZhUPpEqedsLFZm/u8TpeuDtynss7ZG1fInTxjH37Xj58JSAxdpk8L1Pw3xWPtK1oUzmkdwuXF0c
tTAfjOvRdPB3pF8R0ATBNBSQ3pVyUMwlGF2TcU7X0bD6yi9Mf2oi7CqnhGa9QmRRmT4UfZaMELTu
ViPRyOnBuYqeFRvl55oUchw8IRICjE1+53shOMfrz+BmtXYqCwqSo1VYsFS1zCBdgl7D6LfgkuKn
VxqAR5ImoHDhMEYUQacd6G/KMjNL1ZMNhkc1yoI8CXVl/ytnVZKnWKkfyxeP+UziXHg2OHNeSVP0
nvmINw3WT1ZmM6HfV3HNs7s79PULQSFgM4qjIRpbQNzy/LzSpwjh9GMGdImSsonUdGrfJX64++lU
oMuaEh+ty9htrAMavSMdEenuO60+7FGNl9vfuuUw6Vgt9e9IIYb6sSNpwZGHFvbjY1NoLyIHjFQ9
lwPZIQtC/7W8mO8UQxFlatPk/u7xLspvQ19HM/ES7+krg9ti69n0R14ev70Jn+NY7jXg+nE18VnD
0M39ZhHauI4zkcxqeGvUXeerC8xI3hrRVPMVcXHYakFaL1M5x7uDprjYWNx6WP//Y92w1lquhynS
bofqikoGhLVIGpeJQs11mro3qSsJJLcHFJ4EJAAGPAnjSzWwcIcS9Ds7EhqrSj2L9r+nAr/lN5KK
UyTjY/AwuFXVll/Up9cYGkUL+ViSnb0/BqBEkDnLuP2h9DhZqPIr3Z2YCfZS3eO2/lEeKZEfX9eJ
muUwJf4O0lFLKtPknXgkM7Kbj2ZNpVtNtJ/mux0q9U0WmFNLskUgSYKWRRsvIvZeKV5hcGnMl3is
w3xfd8MLjpiKu4pKt4o2X/L1wZKO2rdBM13mK12ejKHcPX3iqxAqGknQqUtVgvNe4thHOCfEjDay
y/xqzQKinAKBIcwScE1RpUIGfcGu1Z23aY8PcZobO+XUn3FNaRlyVwaoSDJWTur5skw1uIT12xKY
ayuCBYJJm4Nwgr8CV0d549sgaI5fkMqxNgJuzX48VflkSUnWB03OirEEzhm0L4sq1IZeSTZQmx+a
XR+gMmlyOqqQOkcPe+QUuop65O2Oa1PhFcOXiRlXWHc1zb4Qqc0cnunEqJ0vHO73OaCY5G8KbcUv
GDs4tEuvb0vk9Qobm7TZ50qScx0sr3EPQM5mlI0NbObbSiw7NF9OFYBhQee0X39FCZaZegoBfc6A
CgUfijyxBH4ew/BZi03cHR2HdVj/8CGDFvLGCi68ngSGiaCnozsvOciAKmypeLiAxrv/ct+NLGzJ
tUL/2VKiN8OF2IYftoPJ5PzU4fJ0V6ABYugRgEofmMTJLaMDFcoAjhmzaDeB6OUbePIF1Wi6bPmF
io1RFuknb0zDUCqItMlOgxU4CD4NjqMwXd2DO7o4GQGVz7Q2uSqJnUlxP7jKdHfJnjhNOA7gfv0r
rLV2DWVcGnTH2Md/hmekYOcuxZ+ZuYFNjlYAm/lrVi8vT7Mv1boQAsz9opTO/CosoVsJ1bsy7U0v
zJz6DOBW79EdTurTNLm6EcaFuvgnNogdsRM02JVZlz7cl306wxdGIs5RbeCBIjHY4+ptb0KpGnzU
MUN+nGJNlmBZ9h2gdZM7KwfIf9Ks2/cW0ogCRW4NTmiUofamjO5dYuoniGm/FdmJwsUF5s79xwBZ
rYv8qj+a/iCrptGhR2c0o2LfD/hBlVTtDr824zXogIjY8ZJL4A7M86LNHWLH4nIEft1FROkfaG/U
FCzm5AxIfd7/5x0cCr7GY42Ita8TaMmMEYZr6Gj+nDG6tuKioVU6NjupWlvyLxFXrrXmB1Uz2z3B
cwevUMjI9UlfLR5KDBwSVwxrOlEuluFD2j2au4zXXxY3E+i+YgAwwcp1qcaHvEOA/Tf8NKV42JgK
WgJkvQfkdVl6fbHn1d21vmQi8DtyskeyJ0EAF1ZsossDaP+uwq2Ni6T1afymYWGo6CMNUyIe4VDl
lxXQg4Wl+sYmtJ0fVcDZMoaakWE8UGw8Y6Ar9h4zqHxcNqRFDf0NctdG7o0Jg3g/OHlucdUr+DMM
YOvIUFD6U4N1IDCPOuu+PeTArLkAu8wCEn9MiJuUaHPmHO96dpmUhm3T/Gg6EpdPoTuDaJ4lg4XH
9QrFydhCkUZf2JD41OzxiU05j3QzmgjANycHiXDMzXmPtppQsCwKdKXlmlM1KRGundlhzVUx4w46
q5i/dIY5Ih+5aN7ttfhyA48nypJBE2r/vaI0Ueiu11egD40tSB3fKOCfKQ+A69pwtJcXUXjH83ti
OwaydMsSoYJGeti/6RIFungOAzA6v35i3axgJwLRlmLQNnBcdzWBb5FYBWqsIRzaZmLqC/cYLyaJ
P+R4dzIh57xhfZqQAX6ge8+H1kga/85fKNBaN45XpVnTBLEgnhmR9JTkeaqIdwvMAht/HRfWRg0/
HEdd2zrq+eGfLHlLRWXwllJmSsCyVxXGoWUbIryXPyKec5f/MDv3uYTpgO4CyHpGOYHRBkPAqMFu
it+9u48MYPVnpHxOsflnSrkd7Xx16SpQHOZtSn9Hvdp1tBLGZbH9khNlwCgijQOG+9mN3bIdZvJz
53iSFP0zvCC44I1IvxYwYVmzoiWM5/0J28ZfMkKx8ABowCeC6934c3TG72bB7TrQzyqkeMaUIFF9
qaFF1JEAuqTeD4QYIH1YUbpUw+gGabEaNwoYsLg7mbgJOpRWNW4+VEUhaDIiwC9RCU+nclikgqdj
jwaaCDMaOQ21rmPkiNOzTbF03XtJbpyRjWtLsBpK/l2E6VGWtHqhEkF3oEf9eeNg1OhWkI1MjfFY
7lubfirWB1jSsKZ993GJlLbbGzYI8UwzA1OKUyG/zB8/H7RowF4mNoQ2B27DMGs2rrWbraFd8fbK
nDM64lJ10IL8jOsPfynELJYGAQlE4lu0nafZoQLa+w6dMtABT6RQNa8Fm/001gMTKQpzIw9o7QoY
9GQ4H5HhKSIiIKXeFxpKy+EE5HZlscenfgyi4tMyWsh+hbsqjX7V4ZBS9zYdQnU2TeiL5ToXraQv
hqCFUt0u3NAfZxPBdyv+7dfzMx0N4zlQCPqeWbnUP+6rKz+aCYFgQT2bzmm8WylEAjbBwcsPCLC3
kun5Ll6eEAOexjGnlfoYpECI9aIEG8rPyPouEoX6tXeu9VT7v/tarlX3fYtu/+KlQ4ayMN9jrf5V
+6w1rnBR4tEAR8GcZq+PquBK5pD3/NBTWfivBxV7p5M5r2jQE6NjGaRtvuwX1c4kWE/4JPkki0ng
K7DCjbiWyypubR6PpgpSOSOmv8439glHd+4C+51hQ77xorrMIPqeIuhjebEdJ5qSuImGu2i68Vuz
6Q2kHGttHIW7zm+X1H5AVcbUOtPoFnU+mV4f86N8QS0hgCXLxaIRudesor+n6GCQ0Ox5UKvI/t8K
isAvBaZbKoMhRsjNWwQr7sO5cLyn59g/HK616aFl9Jfz67JzVZU9W4WYjOB8dMgKM6wx09b4uR82
LJGnClFCLidI2DGSx7dkP15J3mS4D0X8tO9ch66ZKxtQIatqqTrIW69IUpAfwwOjYBMbdoOpajJg
Kai8eETGS7mvT/urz/UFsRlWRbocBGWhws1/vxi2OVHl//JuU6XXTjXbP7R2Kgu1Ty10DbNpx6Ln
D0BYzw9W9DvJZNO1IM5I6X0BewxCCarOm3NZwjiyjwYwIWIXe/kBW7zyQQRo7XOUpJqT6mHShfuM
dVVP2hk5oIxXq0yr7gujA9ka8dbKVczHGnc6zzT24JLnRA7Iyr7VD4KFBeaK+SeX5Delad8aKbuu
Gm21Ydx24ZbidDvF78YzQR68LuQvNsRn+netKnvxU/QtzZ+brEBVOw12ubFFbzOEcAXc6F2e0/tC
L0qy+bLtgW38Skq7qP5uWbEQZTPsdprwqbu+a0UF1L2izvvHYTN2egn0b9LB8oURxw/JXaYFfpUC
olkefJw2UxbohMip//b00kGy4DI68J0IRk87IvXBIqUI3UEV6reCobalIq8Y2P0SymdHdQo6EnRW
3m3m9AQ9aJKLDUNhPvMeFFt99p8Slo7tb9uXrsiJgYAWbPmTjgQt4EUjTqLvl/6DDUWGynaedVVR
gmX7/3y9j6yYsBQr6uTWRssNPl/DDxWKtQxIJtQwxlLyB9Lf362ijNa4XfWYBLMs+0ZtcDkw8Cvd
PYxH5wZFtXuJzh3qW2bzu76DF2t/HrbhUBobMqjPr4oDZ6kWz+8/ZTUEDgLYixTAxSu+jVJMJ3od
/j657bXY7h7wX6UHJpttk5QX+5f2sB2+gQi5dqWd0LXoboq/BtS4oEZPkTRMdImoSL2tWc3NjVIE
9slAfqgquz343I88DhUh/xNzYZSzE0TdhTlwZoXMItbxcDrhPBjzG4F3/1e0pWXIb67mTMKCHalA
2lh52mFT2fFaCceDcUYHyCl07LAPpnMlmjJkllNf+YJLSO/2prtT2e/q2zHfN74X7esadtpNDbiw
fBjObCclocVrUAloQtj/bAZYRDym+ztaX1cfoadHSvOYQ2Ws30rGgcvHIIxiTcV8e/SOlIH+3+dt
yU+V8XVnlFcN0Pvs4oy1CpWWNSPfVQ8tJOfGXK/lbw2ybUndWBi/zSkZVvsmbpD4a8v2j7jAk/iF
ObJOZCX3h/sRkVzRewugn3D+lZYxhjxi6b6LDUBbl/NIGSOoBgHAH2nCJywXW5CZ0KHWZ4UHu5hP
iR00pFfyRrACRGaUaES1o8pw/gBkQ1krX9lI2GQilzgGeiKlJzhZgYs3blGJOY1ZpTORbYhtotgZ
Ccjyg90Sw9hllhq23vIjUsijGwKcRQrs19g3wSgPt0GEvz1kD8MzD0Yr3aYgaFluyK64hYyfBnJX
f6nY28Ijela6MABrIiBXS+SLhsxS72/U79x/n+KRkB6EOid36BOjHjsttYCSzZgPske29JPW8J00
u/NMjLbqbSWz8Ba3b1fGeIz9TSZzkVnxdyux9vBcQmxUWACbml1H7muuaI7Weuo/ZQDweV8W98x8
Q8ldpJ5AV+rqK1egcF5B++VPDQ4P7Ffz7Fj5hkUQacoxWKNQFztSp/MCgWYS2GdbUlfHxaiFGsHB
OVfrNutdX6CSSLuLaVax3AdYnSOpiMaPjLL13PqtkLjUW1KrHDMGuUI6sj3RAy3MNIwy/faSyAX5
oooCwQg2WLTt3NI2yWYENDRJ2UjIs35LSO2qGqMJXkgaNhwG9qbVI3g2K3rNx4de8CN8brvdZqFI
KdoNkiSDFIVjhmZB5ILdfBEV6yzUz1UaIqTY7Uoq5n3lpfa3c5PbZb52FfPU9unFy2TSxYDmLI5+
/7ymWkYhKXKd5TEHJwR8WX30LZyhF6+OcIDsOt1lsprArtHQzE3I6PGNSeUrE72Ol9hiGDjAyjQv
VPgMF4dQ51eDmvX02eyVZp5hlkGO2jXyqOSYZSra2OwLUgXVnlbIkE4wsqbM0pq8PYXiKI8ejZvh
5wSSIyV6QBsIxsO+NpLI9px7bK/Nf5zkvsUi1liTLNKXQ45BFfvzI0ldeGSmG11pRwZ2yD0ucv5X
T08NWijhqK+tzQjb7E0TwZd0u2JAaOFphfNBg0vik+1KOc0jQgR/qIg7uQBHG+l2XKOOroHAyTDH
uHZinBYaUXA+jJnmWSkRK8LU1BrC0sI80eC+eYzrmZxiyGKyn2rxMoPAiC/+/pc/8rJcBNoDPLrx
8bgHzwMrE2keyntGLN1KuAW5rg4pN9Wa4Vuc5rnefA16ME5IGtNlFCGz08wX+bC0RckaH1be8l3E
jNMbSvZNYGcqyOm0EfkW2ZulR+8nvdOxh/ADwCYldqwteaN/fK0fMb0urP2WfdF3j+u7lrseOyga
ztWrzYgCiM+vZsgj9oQw/EfB5fieB79dxcVJ4yBpiL+hmqhQi9RJ2APXBgRUvdqUlsCGCfZc0Gqs
Op4Wv//pUvTbAv1NJmiqwsdj7MsLjMWSBks72cT0HDlSnun67iXLQ39gMiAyEk1F+YUltLPVDNrJ
W2ALJacMYt2FUe9rsQnn8nyW1rlkLX+uV4Fos47BMZ9ZuhbHlv+xRHpMFo8cPzv4kMI34UBWRwb+
U//nPrpCiTCdt7GqmztIjJOQdX6fQwkQDRK9QL5BBIcwoSpuDRzBGCnR3kbm31igcpAEMY5pTgoH
6FZnINYarQYQVV8rGqL0eRL+uVCf+YOmhWT01SNOM6l6baU1/e5SHDM9DP0EYeMrrsxguNWKWdML
QVqYIeKOD0YFvE49SmD7L76hX4O6Gxhra+Hg4qab73TbVOHnCH1PtipQSTMI6qI8j4wKAL9ZTJxm
0RqLmDiXAB2haWz2sKbwZIndu4NPGgmVQlywvykCBJlaOMQ5gv9XVcDRVGOYiXv2gk+CyQpra1vk
i2wMaMAm26Gin9i1EHifWUSkHd1Bw63672f30p/OWC4ifKIPuHV602paYezNYtT5zxtVBehZXnsQ
tQ4/rgEfUpt9GTmyQtkBPMuMrouBigS+zZBjqU+jNUwh4xPjXWRNTADzdz78/qk4rcUeZu4CTuDQ
DBfRN9XHnebPyJE8//BoEM1/UWVuCLTQw7epjkEQjgiAAILqcsz9sOze86ps5skgOAW+llLVXK/d
WVlxFJ5+4rhYu5B61GgXdJXwLhDn+cR2rkUUJfxITRNmrnlKEMTmKIutEqD23LTrfEZXDIn07rsJ
lpkkrg7g1dNmX4ROEV3vJjdnYEup1ZDdTQ6swgYNKQlfJ4QUnrVIxhdy7CGkyewMQIUIJVSzN5nG
zBlGC/YHHeIQJmLN//v7FXZLvXD4A0Ipavj7RkZQMgntZ48Rw6LUZVEPDqU/dynrS+VwNs459KOD
Qa9BPYH9HgsicE67px1+eHZk0uY5A+Fq+6HRL2Mm64viwkfz0nj4yWelZB4ijrcA85QZWxzIx5ME
0Ggmsaw7Xh/5AqgbJW/quIlm48CUpYS1QnMNUfnIFM8dff9K9Ucqc7eItux+RCyDHOuWP0GJHNz0
TjMB9tTawaseTwpQBmLLX4HEGQ5ve0XhieXBml55xjOj2V6UcNZRCa0rNuHipxslFeYkSXJ8XBh2
oEZCMf00rHNsPEKYm0KIXt9fPg0OttgRyQdkTO2KhHhnHMCgA96h9WkGnb1WEWDCLlDScyybxOU+
nzn3PlbzywkOojSRLmWfu9+x47w4mhZhV+VGNe4CccbWUI9yd15W0vDzMbngfS9QoGuxeq8EhGEC
x17p2+Kb7YY+bla0hLjypY0mqcIVGxvPDB4g214L+SQg3W/xR737CNCvfETQaFlPRjExYUf1GXzH
PxTTCSghzPZLE8MGqyfe9lTZ37UdePjb6OghysbsEHr0uTfbrlwt2StWIl2FVbjfpCE+2CXcSZEr
lld/dsnqep0OeMyZcxvI8lj2zA+h6PtFbxtYnt33/6p2nEDlRE65ib5YNVtGCIET1FGwryxHeAct
oa8ECLIg81V/lNNOiSTFdfW4YslHTLHp/fioUikNWZqidopQemr850eSmHdiawZKWRlbqFLCbmmG
7AxS2ZEUGZZk/jltre91JqLkMfheJuuGHfIKAX4gDCnGSJl+ANoBTtKq8tF3y9/0WVjInqbbRM3Y
O3kJ8VeVV921doRErxVfVeZ+7Z1kEmCTA97lVwfQF2/PRDDnHBoFGK8oG3nKEY355UxRtLV4qDSF
lq/+3IhscmzYtITduOqSsbV3B3QwIS3qhfMAoqFiBAwqqLfccfpb4zrm3jthazUWNVUbxqB1373i
NlYSh7VCNFzw0TQlt6dSMIqZcXawRQ+e28k/96Dyzbz67s6m7vfstDGeoyYokIR82YaKeMosTQ51
oFb5UOVHY3FnEkOP0riA5bNIFxRh94UT0NmT59qI6587c2BhN7rDHy/P7vgQlmlHXWgsNinNgNR4
SN/de1bzAwrwtmk+XbcxSbrdlWCNAV23Q8XDEimtdFmz5YLepXx+ORjoPpK1d6RtqTIlFnFqWF+k
S5/wMzdq7ijidW9l01f4pJ6Udn3KxrtdNURl1P1XIopaDU37LpHBf36WO3I48jsGDoYt4eCDTzbG
peEu4WwFNyLsO/JyUyEmBBbr1N0qKGX+JpSnczoCYeInBAB095vYsPhIiPX0nf+oWfbRjhPbmZfT
GvFZMJi5sWY45u/KWglUregx58N5rfvsVOUx5JEH5sWhPQBGF+WiCq8tF/nGXSP0/k7OGjzZDDfN
gINmFGoGyQpi2HJNDcYRooUCJVdpLNYaPomxeU+2KW88sQL4Xn5LTAOu0kWoSOFvr94H7YnJPfjH
RLRBaPsbz/rGwaxpLHs6wMnoIl7t2OVKbA2kgYOX0fFMGd0lPVZsbJivN+HhaUB7k871Q/E4s7xi
qMHY+qi/u0Hay3J76Zgr2TaqiT+9vsekRpyEutA7GpoaYk0zQn7Wtxq2SLQLcujPQOe3D3vqFAAp
twKzOgWegemlkVGmIm+DuVMUc39m1OgtLh4aUwWpdYmWatbTC9PIQpUhMIRUVmefzud9A9u4CAY3
x0xntopFzNS8gt9o71OGedRpdu9aJG8T6DF4CTVXkvTZME/18fl258FuxD7rwfKKi42snFasMN+L
L5RCY0DqA0DHdfYP5yw3UFlJNOtB71nKWzyEAw7FJN37EjlIMru1vweuZJ4N43NjGlGr7Rj86qGp
B01jgSZQ4AOydFg2WaZw2KY2HGTBzhu5NZC4qqYsyxcapPnXXL8F6H7OmQfWHv/hIJQl9FcahoYi
xhlIlCbi4Gayf3eCgIzA1hhgM/hHyZBq3psrSZejwS8gFfh0nKQuGcbbTpKuwhDctQRKtQ8IjK5a
owohpgAMcyw5nKSP+6o6557GblLLi2dxopdL2IB6qEsfHbAbHc7dpa88SgoGRE8UsKqqyDXREoUl
QG/t7KCCaDokGvr1FPBCQregdkpy7ODwpvUJMJNV6tmweZoGhU0KJlxCwjV15MeBmRpk0ql0h19R
lr9jYBYCr8kyXgA5OKYFOdYhDh4CirCvH1xE1wjgHDQ0CcqtLn2qZJrtWkLcHpeE1OFG57xjnN6H
hjwZqvBjmQxfOxi2KSinpv8Ye6rIsr3HPzgyR6nb5jVDxJ5vpK3WiVf5j50GuyMb4Y3G3Dhg3p4b
1nkzL2u+IjWvoiox6OpQ3Y5ng/Tu/aRX+xcFy+MOxMik8jLjZmhpATfgoc+jf66FRyV+gs6PafEh
/DhKHgzvV+ssPt6zdSa5NW9qG5zIUr6tDyDr0U2CO7EqR/ZuxC9uD2mx2d1LIn3bzBKgODZe12e8
Mqjv+w19md8CDdcMWDE/gbEqAi1JmvFJG3mNMW3lZxOFz54krXUtwPSBaQ6O2J+DFdEiAV7ryNT0
BWFZGwCXUAI2y6650ucNKVX+3PnY+X4X6FPOt8M/pvqgNXKh2GsVQ8F5qdKue+CbUvJfXlGN+rs+
18ziLtT/+Evm0/e43z3v1wjinFE31AurPlTJrqe79gBvKsCJzzU6q8/tN3mU2bqRvEYzO+5vLneK
bCNeO4DOifuz8x5Ar/kUG0jXje0Ca41gLWKoRSpqgxGKctwqKsPl7lTUGeCc0Go0npHRj/bdHDoE
rsoAQQ0BEIikvDimziJI1BYcjFDAf1cKVYoi+k2oDZFssCu7ghUVidMlEheFjPka41/r3DCf++hR
XxoqTjKNHRnAKnd8QoOmnRCnep2aKKUC8xktigoZKW+FKigMiq6U9PjE0gBgeO1nLhcxhCs5NNLd
EaGRP/5UTkq0O3un6dhU4OBsMNLuPxsb4102kmOc3HkgO5pSDTAoR16Z4MhI3DcTfMfGeNeY/wyV
ksDZ5sG1JWIrP9UtkUpHRFM4PJ6a01Sl/UMUkp/wE45QyzqB/iJqk1sM44xVOnZnMVgxv94RBLix
6v8xv3eTMFAvn56gEPU0CWNodAoQble2pfaLzOGEnLdZ/eX36+k8T5Los/8kKaRzpzstUHPmhdV8
iD8WQPiwhEiRYBmDgGATqQ+ectH5gel7J/XCuek3fBkQi/xFypSL0JKFsmq8tw7WL3n+d3U6eeUw
9YxQoDYYZiMdP6lX/DsshT7M38IZsTdn3RxOiQwQusHdKRH5y1dMJRlazIDpUnwCI7jOqIZc9nYd
Em5BfS9N3irxbi+htIANCNN4y2U6q1I3WQYuQgHhQZLllHa0GxHY4l0pNp1o40Ux4x79swaN5LHk
sZWnOqbaLi8WUqzrZLu62aYHtd+HRsPLdi8HJ14NbcflWo38wGv5gNPFjuKfVVio/eZs734Q3ZDu
yDbqzaP3LgrkZLYGAhWvZpESqN/KTM6ZbbF1507cbDGsClxFqTV0LSz/hMHAOnJhC7hDmykWkQuw
uXf7Tk4F/jCNP//CDMcwGCoNjC/REMD2kqw6DeHbYF+zvXhgH3c+M1Rc5jjS/LYG3V4tKBrfwGCU
x+3jlUeM8oYXyGcrEVTWsRPtq77Dgt3/PXkRMHDA+BHSfqVQDnipLmnO98oYLXg/Nt0hMt3Kwe4N
WsT8z/2ajtQglk9gNH/T8KqInEHtFVcbu/DqbpwWOTeO2FmqgB+Ny+IgaIf6JUOGk8GZEledj0LU
UnfGikJIFfavdrSqcj1WfpDMzYuy0W0jZiE6YOGgw1Jmh12dvcLUd5ZAXFh7MW3n2joGAEYYBKf+
pvtTgnDparlyQylMs+9d+mqkLEc+XJG1J0NC0e04L6iJNMqbTfddvDjkpCzePXc6W4nGA//2KZZ/
i23yyh0cbGufJ9s4PbHC4VWaYU6IRJ1rHg9avNqEGdzgxniWKRBP/OIe2Sz8ijWVZaoK8e8PtvPm
RQPoVXjfuQkkPbOcarr28kWK5C6pKcc/z1RTQ4UD0EeUpxXsDLWJbbXH4Vq9ssBLoeU5PfPYiL4N
pmuuedYyfD/Mo0hKU5LSAlYd7WZTc3MCizeheqHTLBKtOHAUQPeZecDyrjZo96SYANvYyci41lGY
8TaWkBwo43K5YErXtNC1GK4XJ5bSxtBqqS8yaaoPVazkcDEOGEUIiZzkxReM+haCLtRJPW9t+M8q
c/nE1YP2eqkvS4ASo4uaNQguzPAQgMGMaB65Wla1Qbd9VBU4wdtK3Dqn9GNsJTNsxIb7wjEVhfei
0xsPuOPFGISyNakwcGuSNxYqkSUEhuYogtuFVUbkW60VjJC+YXurZsgV9wb8DXrhk7B53fjNHJJx
USt8p47GUhCncHwXRVAPlwAe1Ql8fp2NuKg9nSI4IoVStvzZ0pHiTYAsr4sRB7Dwy8Cy1dyuMXZ6
q9IXfE7pEnIQCz8ZNmShoUCTrcqh0FzmhrIYJMyem2t7H9aml2j/9KARdkojwyBacvBtqE52k1f0
DYyrn0Aqg3oKcfwunLDzyiGkNmo6RXJT6KbrgrVnr/2ts3XYDRLctw3hxcefs0QQ87QCrd8DbVa0
4GxduYMveYdk8VHGIyHWnIMgv0J0XFg5QbQeW72vOyTx6Mnqc0SFbb7F8ZJmS5ZJVUgMS50Z7Ij3
3nAOWKr4BVMlpcBzYvQl+BpvSms7nHmaHMDUpFLj70tj/VDxWTbj2QPulKM3K/r+dhEelIcyOi3P
ynflTz4Vs8U78GiCOVTQxEPyVv47C4d6tKBf3GTW8AI+y7QhimxRZXg0xq3kfvSX4OdT6lVGzQD3
VouPq5GksXsnS4Tmnvuckgq/zH9lhX92h/vcKmyyELhimRhxEY9bPlauL1hMm4ljmLkUgxWYikFz
SMqNLUqgnqktQaNSqF+lq3kI7xZUeaSrT06Lwz01HBjztPw2bQ4siQAhGphsKwmmkaLEhOh/J8we
wYS9v5G1Qd+3osB1RFVVUti/qoOrACBA7tgz9wDIbAZcfs6tXIDb6t6I/DAkamcHeQfjpnbyfvRa
1o6kytLHXZ+cNF7IrTryXitBeYqkaxgDOdYpsceCgqB4PUtPi+ll+jhGzwgzWHOwJfAUgkqWCrUy
Jr9AqjvaRAB4PKGVUI7K4BI7oTyXJ0CZ/j0EcedCIMdoVWsbJG7ZkXI9duPgkBwhVkhrDHMVwt1G
DBuOdek8fMgB6jxrmlYwOHi4jsmQ0LS0BETcRtnh/DTEgj2TnrjPp2fcJ+aOriNEOGTkzyQbWpsd
S7mkpOuG2HSqLUs1OIuLOcdPu1KZcK8iHo5UImWKwqvtAzuHK6+Pn5ONlhx0gVVeSiAYPhPI8pKV
Vs5sGYRc1WiaW7MUkjZHwZVL3mDQZGbeP6dKNrPeX05GEM9I+jsmm/ggI5FPhiL5luPxVnFFpEak
4+LxQPNVV5wT37FDR1hSozTbGg0KbYcriA3NnBiGxYqW6yehXoqOljtxPZUDhHdkIAzOfLIahpKd
ap7gXqWcTukBdr654GJMfTpodk3JPsZg6uA3VxF5gt+k55CKrJI3q+bDUI4EV/AtCnKTqLW1Vo67
vXszW3s93WXCWiHtJ7TnFkHYaWefH4OYISuex6JyHwsv/WfPnA/ztCUAF47Q26aOYwj395kQKi2R
jMb0F70x1YbY+Xnb8rSPnfOoO/vwVWefG7C/1ylgJVoBoQxwVOAOC4ZaJ0mmMr3o9vwisNl6R3k/
2saqMW9+6f8o73zNLLJ1+6lKocml9khKrhO3+6YTXSWEH9B4cGy77HxTXujLd6Nihzx7Hk+TE6ps
8BTTbNyA+nKQ/RUEgw5nYOR9DHxViwgpxABBuQxaYQM1FbSWfsajXn1HQPGW23Lzd4OtPPWvoJ2b
pD/0Yj+QcrE29DSnQhmySlvnJtFj5x20GrsL4KBt/7cHFc7U3M/dY3n2R1Gw0My5RTuUJHXcqfk0
x50TGtieO8EEMwYe0tI3t2f81O2wrRKUJvNptsC4YOYP2vy8ll2MJrNIP9PZCd+Y0Co5T4YkgSas
Ta/Di/vs+nLr1R1EttVAAYdR+HqSbnzh7AAn0Fb/ZsuhJ34sN0aiBglGefae1eUhZXz55ergZS9H
SO71KYKack52hrjcdWcY38GgvjjoxV96jAWnEdUi6qGLXAZmzQ5xtBOD+AQhFcDuEoySiWw+8Qne
+B9J/g09waMbfhalHeaLTayrJCRbmyIxU0Nce+THNQ1iOfn6dK7dG4QPyT/l7/w7/gR2ZXNL5HsW
jOe1qF/06OFV8K6XVaoWtUK47gdGdYlk/6fA47sqFlQLIZhq9PQPipcjoDaFH3+boJifQAVvmvzW
vd6W9lmUZH6jlCbuJxfE4Up/8UBFLfhycU8xyna8MIlOVqhyO0uZX3whbrBl1lhfK8/ButA3lQjU
+bhRZ0x0AVp+Jx7QlWzVIj9hr53C7pVK887Mky2mzD+TVY8kj4Gp775lnWSfBwMIFnh8Jxl2vVpq
e8KotDiyVKDUk8udvT09osZhTnvUZqh1BmX0qc0dIGOBNvoyLHJdrUUrcp9wQ/DIKpRTc5oOZJkS
9QdpMSnEVbalH7xg7VZvlAe9KIWPmn+80JAJhoSBKSs+dXu9eJVU/95dUPvpX9jiHFilV4ZvSWx9
taRfnuLa3oqccmLw4Ulih93RHmjT+BiJdNPZ2I2Am6V0U/KultLFZLpH0IENI0twYxK4HB2valAo
Pq8Ngk5AdxlQNQvHwD+tSSHE+Vb0uh8pM9VusM40sjnD4YMtA5xNzRDoi92r8chIyg0UTycPHrJD
RP0x/UQRdGctwr2968UnfLT29cfFbeNsj+nRXyok9s2n+RblcT3rHL3BFBAnQdoaLL+lfZimh7Xh
pjlkTqwyNtA7FVJaoLPsK6weedmBsRky1d8Tm7Q2YLDgYaLRIOE9m7lfVdqxuEVUdvCvLhym1cPV
x9goA2eQvi63CXN04kvVr9Zc07X5gmibAsHZGDqy0oh6y6lMv/WGENRqmOTba2kKR26wTli9jaIB
m66MRNdz7Ao5O/bvBg2x7KzKur5+T1+15PBUWb5ANhbTIdkUZDMH/n4vOle9ia5R7wlI0lnDVgYy
5oMsKNH7rN84hHR+5wScHTf+/uK/4Vwj58qEBYb/TqUy97ySbQB/OPmQiHeCPPimFtPwn3jd8ZnD
kROXfZXbndkGWjfq7WiL7DPFG9iYXtPE5ETDHs8lxeKOL2IGeQTzICxIFTlOnxmookkgklpCk6+X
Qwmz3LvXElm1J7u91owaHdg0D/Kpwq1BpXMbVi4wTroNCVJFg2/eOQd1pewBWuSgExVQP1QET4p0
HU3hNL65RdmOQzDdsaYikslw3buak+8PcJSdJOlb8xT7aQRWo60l6vvfBj19OB4AfrsVCyIfKA7e
0OcKG0M/12p0KGqdg8In1CxvTP6ulQO8fnfgbsJ8KeotPGQ2Bjo9j6k0bG23pqUIH9YA7AFA9821
o2nytNgcH3/SNCCk5bOybIbCmMSdrcvjsCEjzfzIyd7MD3ORSyfi0ep9KTJsJhR2bFUef8WuOpQ2
mrY2VdsiT/ZfgfGuUoJ1qfnGcfw+e+MDO89V1tEGadBRfo1OFfpHhLDpm1TZjz9Upd1BIc4WoMpP
NHhy5b9eirum3iwuEXteQryMWH6QqzYPausp3806qvD5bswl7cTIZqRzC7J/sTyjFczGTb2ZtlS0
Cs1BXsVWvdp3+FB5H+ydeEm7qcoGH/NSdMfa3C8Rh7bEx2weVhAUC4+LPohDSnK5C/sGPZ2Bc4yr
jilo6LQKpwgemNsesXCj6R7dqhjlWXUjomKyVGNnZL2BgLyOwPRwakImUDiijTFg6VECkCI4hNe9
gnE/ejV6128laezV8/hpy3Atc+oxBbvSXwxYHf+mxUQljOrbgvAsJaKlGYXYwYp6KxlNx8WjteDX
nv1QIJA9l2k4mqGPyfAi+lQBOLbpKQ+FqFFAsps7DfW8/BiVzE37YNzDUiFCP7rarVlar27ehw9h
5ldhHLbeacpd1E9YV73q4WpEfdPbcXNfvpznKNdbii6IdvoVr3VPCcZoN/L3H2h0Xq/3NaztETtZ
OS//jccO2c+DF6rS7G/3U+dSekZnyLmG+4OwG6MBNOfbOuZttxbP6p9VFEufEjsL6z4UD92wcUxp
nZR8hNhHxJj0pjSfHfnS+Zr3z1oV2JlEBtQLGibnrQWxUCfc6vdK43MZKQ4G+K+pkOuG8laMaCsz
qo2SLs/154gpXnb1wQzU/J2PXbvxYsijpNjM3GwniTcwtN7B4XIJZQTz0m5XKtc3X9ouTMC9ggN9
L0tmHUXtHEiJ7HYVDG2xIZY0Lp7BpCw66a0s2b9nYq6TrAGmr+VU8NdJRBr33r5HRF6zQ/hD8QUB
LwIM4idQLnDMeHWRwQdi6bZ3IUuIBVUUhbBiRtnWarmKY8m4cM3K4gHLz2dn8kBQDXCKhwxJZM7X
J8y3NJ9+cae75E5Fr+s3nGwFujYUKyWJCqVyEullgykp/WFOKpZgFW8apl44cD5omwNlmr12NXcs
PZXJcqstKkiX91TFm9/XEHQAxwmf0TxUFq2hGsBrYIdNJZ3RnyRJRru/3suTiW3xqKbv4xRSI5aD
W0Re97uBRGuumnep61nUzV9858TrZpy9eIQ5jLSA0NqahcQe34hciKxXX+PAPd9p2Zp+kNj8y/dI
03rheX87IddZco9WcaH3TGY3q0vKQ6iBSiudT68oIVqkckxJIQX8JG1uOCqM6JSgW+SMUxd4eCLg
DqqXxj0nYLGyUiDjj3z3c8ANiLAQum2DMmhyVRw7N8DvRSwOT3IDiZM6CuE8PsDdIc2a8OiY0hVG
nC3v/CgAGesKWDbu3hT4qMfS7FwMMCGlCfoBIWo2Qb+XfEK7eT628N85dCf0DpcZ0qgUFrEeXJUX
q2+wO4UE0+G34PPc8xKFVg8X0/IR4Z2wp+k5vpsJ8atR41dEH7Oi6EMXlKMVbFa78myP1Sdwr3m+
DdP55fh87byv+dQAC+pEBVBe8Y7srOWmTdPU73HceeHJwdqlJYTvUyQUJBH5rK2N/a7+IQPfj4y4
0dX1auaAhtl1/BdHd7GCnvkMw+Ny9+0Fuh+0MPJp/aYRSjXP+8skGJrciIER3Gwo8sgi4rEac7Ut
zz2LQi1q9bx7QF8kuHqYoVwGhFwPE5EuZzANY1Osb26wuwphhhrplTdp831e94canra8QfyXPglq
ViNIJbnoUucMKq1Lk29VX16sqKvod30YMOxg40ljEm1BeRjVSfizUWaUYq0nZkR1aOuowTsPBSFV
+fOUEP5nxwqbwmHfBto5YzRBxNb4vLuEpDNih7k8YWoJRSrjUJ+LUmhbb6/h4JRekytoO8u0iSfG
4xGRgwS1Wn/bTaqEvLR0byVUH4j4MkM9IA+ugGoWrZEFlGc0PTRhBQCzNP56dnI234XvCMTK+j3i
h3iLUxmWdIiR2JOC6wjCii71rFoAsTyegt1hYWMhQScJG7cALDNVsRhGI03vEqQkJVslesaMLrCX
cYGhaQjXC29i3Q7Eu1mKiw3Jo717bFitqyUkp3eGoLepGKQPHBuSGGU8fm2GvNDwHiLU5YEyxiK6
uH+PCGxk8YMqz/4AZneaBKLjojYe5PV+DsSTANxpUcULwDS+LUjvZirWZ8AOo45s4OyEw6ZMqkOk
dssFsyqc78IYtI8MNFCU0MxvW8CaAjmVjFS2z2t3JMiNbbVmt9M7cTwJyXXwxUqpTPHw+hwrw1TQ
9Apv18wX9vPtvvuUCoGeH9Jb2WQAW2yjMiWkZaGX27IbyB+oQ2asipDCtGY8fwW7xArJqmG7G2Rf
Om+xsSoE/CMTsNwjzVcfkzLmOR303muEkWbkZBgDWHPvEnFwESoY06I1Tvh2EqfaiPo1y+G1rng0
VrsjbfHyNo3FrlqLFpi0DDPosACxTvEVpQNJ9Cg7P39ZD80snoZaSOeERLIrML5sBXnl32eQFTV1
wnQ3WdV9Ps8gx+LsQ8bruMr/pW6kQX6O6CHo5GWydSaiyBpvfTWdHW5Ty35ExSQ2CLsG6oAusRjF
CDLysGQPviXX4FQiYbRV/i4ZJemScwk9pxQdCUjoT+N6nsV8WGuYALtjtIF74yqgftW1D7aYsrVW
ZinhWFrLFz0R3HGJrYOTQ97+Hg+inbpoLqcS4Q0pb1rUt6yzcjG8GBNCf0bZWpVkPJI3t0isR9bd
0JPCJposP4aDwUGRAFc3xyTem51GsT3vUQjc+2KYdWVpTYCBm0JSaOSx/wtb3IkR0aBGHokRStpG
Zrns/ZQ7K+TV5nfOez9h0oAl9lbVqFijLylO+GEUS4LKs3AzMD2fPyy6ZSyvN+2ozXD1S+0uZ4BM
KDS+j46Lb7Qu3mpgZeEImav71ZM4ewDdAdbYeirWpMm0MacTBkveTy50Qieiic5rOP7bk2HH+MFE
/Al5lFCg5rf5wd2TqC4bm30ZNKNfAke4NRbdqu86aRohhCaL0CRSuqmPAZ+BRpiISqnZp5Focrj1
8lQUQxhrm/I14TTnnNx8dlZnU5QczXHeiWdg6fyl7Tm1R1izDTWaJd5aT2T2Cg+kLlW25ZPGnjow
/B0WxckNsLmSukfXU+WZR61jB1H9kdHbc/Nx8maKG85ti0/lImg51qx8qT/ohveK9RILorbQUAYX
g7D6wtHiFSNsbLD29jGbRhNq2SmoWOlOXh1AfCN/MGIq0RAnthdCmf5SQiFHiptQQfFachLFqpAU
wQqSWkpCmxmsBLlprC3O3y1PHYER1MJ0FdxrDI2MBIYSZi7EQKRkjNbI3TggIUscgbYhQpJqn0Xl
4Q3SoaWpt+fzRQpkpbQ8Bqr8Q6H4udyXFSV7Drt4F+rLS5tWHjKROuSeJX2ycbdsuJ3yoq7fj5P1
A6JmdvCByBrH5mLf8vMSuTMRw4O7DabH7eAhR1ZWrdB43qnV/koZwCZYZpZUpOpY5jH9ETohmLi3
QCfrfTtmjf/tN5v6qnufjULhKR4WJW12o8qtk4R31Y/4aICqPRhXLa5hUdnhCk0+XyDQwWecOkNj
2SOtZPCj/E0Lbzpvrjn94r9A/v4Uu1bkBrdQcNSVjAEEeky4PW8l0xzcfZW2aG76YCBSraBc3CLS
yr/sFUUFnUPUBfOrW6d3KUeLQXPNoroTacdhPM4X0XtQsDWAW03SerzcRmMpmSUQq7VZ3o6edNoc
h8W6xH7OSq08qCeWSnLqYQdiV4o12duqgtiV2RsRU8w3z8y0QZQqmES9oZ2x4nuhRs5ngRToRY2D
buOSUF6ExXWyMeoI6jKrYm/J9DkbcYLpEAzbxvuH/zFHUPJVkmae9elpbFEgnrNUEstARoJreA7g
nvFi1h67pHylaTO5WIC5RPpf8YMdG4Y06CfH6IfGwfRrEHfshP+IppzBoiHhRz7O9MK3E/T6N8Do
2FpTEgICT/19/+MsFHgsvUjr1wENW+Y4ssqKhJe7BKEbp982GTsDJrlUHenGZ433xTBh+UESKFLU
HfyZnjHOPyEwsaY1lKfGW+ji/skVPcmuSsfigI8M13VoDnbLL/DHnOsqR7P7NPeHSoXOSuuI+vxB
Dhh9NQnzYpEam7eGn1kfiackSqoq/DUCSY9iKSRsM+IisOG+t2wS4Z0dLPGT0N/PF3OD1FbgmLO2
/kk6bds0LhTFvxgWjdISEQMHfl4jonS/V1FC1dXN+Kp3c5suU8GUQ709IErIxUm4JdCEk50CCqua
45u1vMkdXQpmy3swVHNGo1ySSd7k8JrvOXw9uvq67Afu3BfP+4a4GeeAOEUp0NTHZOg89cbdMGOU
z7UX9BrYA674FpXeSUsr419UgBWrdn8GIp5vp9hT9aPZHea6/SLeSqNsMSyGuOPpR8dEO+iwDzrx
q6FDNmczlCdGRWxiOTyUwBq/kIjWP7dAcbfnWmMMHmpwjEvv/vOolDjPU/QV4HNb0Yn9dLQ649Hj
PGQUhIFXVxVRh/6nziIoIxmMgHVlknII9GblMYoj0nmCljl5ojyiztDFVmMxAQtV0kHprD1D/852
cRYP+KGvBmND8jII+ndFJN31enHFrcjMExXbuOOSQ+H/RDPw9L6+UAYgthBycOtp5GQqbQmvirB+
qRAGqR9RTPG4APa0ioUDMO0wkPFZJQY/Q3o7NUKudkNEbeeElP08KettX3ptouh9yoRmCurJWt6k
vQefNFmx4xBb+jwNlyowU9fGXz6/+YWz+gE6HThQe2vkB1DzOWwJ8ve22rDC+UMij0AchfREjrUe
wk9Rcuw4UR4hjHEYK7DZYWz5xpcG1sfoGwwusMN8h+0LZbmvT3cozR9EzIq8vfw8eBuCceM1M2TR
B52ieXk/8cexf0ky9xF1iRIU2H3Rw4EycMa3rz8tkkpEa7Xa0Hc+5tptStwUBQmSapuS4jPV3CIH
qGrgN2pJdGon5RsEq5B6eEJUbgVGcdc0XS1CitcVI5Bubwd3NlG5vRyfEOsRlZ0m9GShQ/fazLaF
rbf34/6NuXGreIAxf5VP4t4Jf755GIUAjEn5Es+rkAoZaff5N4j9NYo+QoZOhoFBLBanSgXA9B09
jQkEsjlAZNbMWIOGHbr3ZWdbtyd2CibqN1HgXuO3lANpOOul8MejQ9P/kLK2ywHyGtROyxcT28HD
/v1O8i/zrQRFtmzhaZme2SDyAqI9yDCsufsJlKD42HGpS1nhf9J+isT0IZFLaUp1SQpADKc5rnUi
qxDIBqGku/Wrv0XRbiurBIrkExO2FPVxWdRCERrn1ffNZwgvoaLEaabthtpkR+e9xal1/2SjaLrh
iYQ/ytaWzP5rByRbvBBrM1M5bfdaGHr7Mm8COnHaCl3GijoeXZbOajS39JgIDc9Rv/bU8cOyEtmR
LGHj+0loaS/pn5CDS7qost+7dQjNjRpTvertmBI0TZx4TXP/i/XN9rwd686PW3tLwx8LU25hl57+
lIdIYtu3GSVojCAvHVSvXnE471TFGfJzu4TQ7+atIB9w0/V8BsRS2Upl0ujxBrflww0TmlnzbA5W
3CsbpEVVp1/+Qejp+pNDaAoxa/Dte8TwlljNNDs3UFsH5K2FEYJa2eU9cND4ZANjp2J08XFJxWeP
GPOXCEQuw4A9rJ+97R1GE3w900TNnyHw1wHgVgUQrHl7+GGZBLO5WRrGCQhn5xM8dVrxklGKhHH+
/GUcOS5wEw1rWS4PBAvVSFRFQBXOr+zl6aU6vlogoT0SOovRExVON/HDa85CdDS5mbxlQmabrK0H
pHznnLq3/xo5FtxBEUJcLk7cODldB6Ngu/R2LH9FvSbXxwAxMwFS1h/q1roTxCyedIsXLyD4F9E+
vmp/kwFSzUM6TjE5Ex6inbnIowXymtBCDdshPWvW4gWX2iWvT7CK2MAmF2RwLn1b5riyq9u16rtw
IzjJdOc87BAlSDGAOjWyK7oNrofUzXAXkMmLnKYU19gRhlfqU+Gw8d2mxinJRaRgyN50xYND9Bh0
NkyT93m5nHeQ6PLZKFIOPmf8PJFqPOCEkaW/1Bqacu3lNOaW0TrQ1VWZZ0cRBCb4FB9A0PedI/DB
Mnlnp8xThXec1gqJHi4VVPMKaAnlVf9cZtURK8QXUDPsJfrx4vB0BqOwcdd9DsfmSgJ8OyS+Bify
Ml/rbrYXFHdQ57C/91JNt8oNJWUssP8qLTvzUeCoZC2p6RcWgoBga0Q7BGWn1X6nfGFv167FKQbt
gvLU4ASnQc0aFn9WTaiZC93dOrXm/EGiG+noP03qZ74NQPbfs1wXrw+exx8p5L4CJ6FoKYQUhfQC
h9H91OaZsgUgUXOhnC3Uam+zBLNLN0bbDgVWoEGHBxcrL/KCUezcPEFHWJv9tWVuqXdNBaT6/xjq
yw4kGdkKGwHRJJDLDHYTEQcVkj6ySslc7vnEmwrVwEee2IZWmbwoDiZc1mSGQjB5hS6V+xxPnsq6
yUElTD/R8eKftRb4ycHuuLtS5byyhPYtf3dxEIPLEMnDtT844q8GIYhyvkbrkkoFa9qmfZuMKS6Y
z3nAbHeOEZ3jYve97OGc98+hHjPVVqCO9qOUnpnS7+aM23HnEGatww0kcuZncAel28V7QKn38/xt
ktdRNf7/+TI7NefHuguQYRnk06LCIzbW04XVpL160gtSY1TNFahlgSomCW938H0RpnEt8BC0G4rI
DeAUgGNhyoY4gTjfBPHKAh1N3zppj7sUMzVMcMMkDgZBQJX4/Xgt4gTlveHkjTHrZR2ZfMzgkoqB
RdxhIcdNEJwR3aSDeKS2NwMdchnPZoKtOVfjxCffG+aMwOEJgZjdtwbi9TypmYfzqC00dC9cQDG7
N00A0sCN9DD8BlGAHUMjupzmd9rLAqU/3zc4Q1WhI8sEUTBLHxpabbx8E7d+7KoZ6ULt0+7wA0Dr
4qdJ3/BzD8bMUhUzJyDbZdWUSQxxkr4chMWYQTn3LN92bhwxt5hvLhFvEdnoYoxvavMNZDCld21V
cYY1qeUSPAzNd+mKPZ1ZR9K1Op5ayhdRB+vWvA4g4UfGoXr7uv3/3vvqg/MnZVpY5LzH2y4YnzHx
LvdUAAavlSpwJdQlUwhcDJvpYQl+w+HJ9uWlio3yZduoss9jiUQbNdtNuFFJG2w3nVoBoeuYtrHU
6khCa2W423EA/Hhx+sn3xFNqNW9zTKVJlkq9DR8s8hdf0XCTeJBz1M/z23gjC7C1mKq60rM6aAAF
wT1eDdkJF3v32N+XtMh3EARPATRejnmLRUs6o5hQnBaSHkliOaKabDTPZouiIBgDc8zcZ83rrwTn
jQxarKGd4Hu5xU2F8iRFI8H6DO31Vqieh2yMRjjd4gAAgy1fHd7cOAsY/62jh/QMDVXl4K5cxkHv
KoTrbq0s6aTMlbXy4XJ8c5czCZjaJK/yPmfyT31/qh9U+JH3/lJAx9XhYs1nK1fs5R6OH2Srjp6a
YLjFuAhf1mKPrU8PKjmib8UghENoTi8xSTxWRgqBBA/k8PykAS6R29UnSqFwR8Ke8Ob9/cqHM9GS
PyI0b1ZxaKZhpzYSCLSM/Zs4wa1+a2v1lp9RgGylfqR5VkXPPKxQ49cERNr2K55GXMv6VrzZqyzC
bvhiXE1CDAkz79vOCqO9TueB5t+IfEhxQNKOm5Y9y83sD98QyKoz8vaAZDfHBxn+8I1DGNY6rRYL
/JNordK7khfsmhWJ/kMwaRXnpDUouIp1xxJcvO+X/g3b6a/88J0FnW7E5K6BJo4kTI7hebrf1jnQ
RoSGn1GGziU5UW81A3+RTuaE9PuQ+IL0sEtQfMK9PxV1sORdf146cFLOWhnFoKBoWlU0fprVJm7d
qNz3De+jI6fw3cigHb3HgEg7eIKeCns/Q8hbKQdxUqU7ntt8uaLGsPsYS8aCQUqXyntsRvoKU3/8
41EGWa2DCYF5sJAr9n4lWIP21SSfeRYXHVH1NpjcLNbocCcPfOyBwokdKRki1xfqKXW3UbDy2Us9
zflePdmMXpofDMLnMxAS6hdwgZ8YV5vIXax/DfvUqVVzH0mTmztyyP0InwpoDXRDBLThik4QXt3z
3sycXTHJD6qHQS19tFrjWsZUrOAV4zi5T3llgOLDT4NbkiV0dPWst7zm05YG0fDRQtFynJGAwsiY
gl1HV1s6mK5WNIBfE3Wh4FaiokM8iYgOVXqN3htlW7ba+d4GAtRdTxKR4+HnhmdeuhycQjJ029Le
wT7MMgT0JY6mcW4NoAnMEh09UfQ5w6vW49NXnmGi7nDj8C1QfgmKqzz6adEkcZE+5cAfuY708lwG
p4fob2lQSvi+oGO+Xqf8oUYt25cBpisLAUIcBdEw2Y+aFeBqVpnrqA7Lcur30s7+YX9N2y5H8BGk
WkyH7iUR9xhdM4nfNS+5jMlO0UhxdChV8jrFm2HS2EX1JHN16Z4jiP7qUmnhg69YJNBvC120+5dC
HJQMe/qxcSQgMvFOKj1e2hflLZGNnSzbfbVZpMJE9nbQF8rcyv7WYTKrLz5vcEj+tkVUiCQRY0Sg
zRZ7N2GLPmrgMoUAcWEUKscKmI8cZX8q3WcHXhfHf+KCcq+YkuD6YnqFjHfTqUJhuvpzu+rEcjpP
v0V8L1TIZGYLbF8FIknRgmNf64dMMFzi3/0gdtb2VQnSeBfneN7Bd1T5WlaJGz4rOxCX+jewBI9p
xP/cwY/hrDkpL1bSWd6a9gqAutLyiUxNpP7k2C2ia9clc1MiDJN0saDHUTvkqamImQwpmD3z4X2Q
vPW/jPPhDLC/mJvUy3xR5/URIXcX1qieOugpFE49XKccD5SUG2Mg3NLS19IcP9isaWqS+/UZvtTW
xJTFSuDbYGvLT4jkVuqLpw8v3iVgFWRvoXlYOzSGyQE5/Lft2GJALJqyphkBPl6rpAJaJDBSGj98
jLTWFnmRt9cwrusSDdbmas79VYJyjbOq7sJmCs67hvcNq1Hp46b1gM0J3coOXHy0s43N8LP3PXPd
jDofkrqpnc1W1MtU58SVTvfq6m95t3D2xwVpWx+3N9UU5po+8hE9r8REYwdUHuLt8u8U/ZaVTe1Z
zQJdUZ5PukCkgmMR9xR3BpGRiJ27pPXYqSOMwP+z4tcEnQLV5vbHPE7rU+yGxlr5WLiL0Mxx90FU
O+wsX1CTD3SgdyNkxzAeQ0D75A1Zq3MVY4KFwTsp03VQ9TkVvl4hW9lNXkEGwiZIQ46G1w3RZiz/
DCEwkMBtkUtsexWPT+ClLmwlJ2BCi/1zy16YAo2/ddi3rhqDWjVPzdEKahPHCy/ehNPSC2SEbfFO
imDadTirr7eeyWfn+cJqPqVJUp6kfygNk6Okf18oU6ml2PEPbpRczckUntfMK52K2u1FwtlR2Kgw
6mRBqoEwHqkuN4toaQy6WIVc1MWteZLpFK6xZchkyYOzodoupImZosRlaxH/Ioloagu61uO8UIsl
kGf0D5z229zx1xmZ7NVQaGTRkam7gGUjKSzghot4nWjTCC4Z5AV7jPAhCoVElHTuOt8PIBBNnjxv
FMABIEStA9F3AUl4NeKeuuUkbQ7NnLPjlhfSfVtadxXRbe8t8kpNEbhVwDJuyHIDC5Ai0o9oZWzb
AeC7dDFEWpVATF+lPzi7OSB7sJ9EsqEKJISXawzDAmkBXknuM/4WPARblTKXiwNAjepbrRp+pJAu
K2HkSJcZCIhXuVWZ6MmwMIZwFw3ECUhGvXC5yfgEInyIQpN9VeUtzTkR70gS7hQL+vLKjwq1eGjw
i3u/3+/QCIvaSMh6gE9ruVuXjdSgrBXjdMMjO79vVFBt+94GNCc3+7FLByOy6STXQ8JVXnqw/Wbf
Yz+0JJpiNUOlEvG3khy/zmrDlqpxnGNAObaQfO1A5uzOEMpDuj0jkmbzqrp5SF2R/HMV9G+2G56/
z9aeaWU6YVXrpFjFDGDW8vwdhLxZBLcjxRgnf1KxOmi2YT9mLQcgUbQMeMcO6MbyfyvDkSL1bkGa
if6omGnEpl9FFpLnS7rXk7CqYVL2wLcFmI9herClrskvJhbOCfL2ATW8smsFSWPdc0hhbTaP7ykE
Tnn6mGVcGctGJIbNwOaclbAEewEZowNI2nfsmi7qiVQsUEFEIg0rIOM1Y6THrouz3aK/3O56mLcJ
heim0cnIvsqalPLzOy41UrxJZEZCqy/JIO/gajGneUwyw8xD2nO/KiBrlAWD+VW6yQlT48sSJNWi
QJJt+o4QSdJlg7uMQG5zFD3yOI3/qYOPobOJhSHmmZH1BDNZeZ4EKFu+0ezBPxXD0gQN9KLJbHh7
N1CDxesMrX8xl2/CXDhYPIKZJivrRECctNm9gXTd2BJBO5L54I5JmliPNxwrdjVpScOtZqBWifBw
GivyzDns3CvNRKXG+4mjWZg8ZF85LD1PCzGBxsn1evbLECUqTkBGpGw2pgNKv9bUdo/81/drcFu+
6E4ofY6Indf5afE3yd/M1GcHD18tn+8Smb5QmHFIfL8h5hjZDV28q+pXKS3TqN7GOgW1b3teXig3
D54nHUVtvrkWR11KpHlzcs4cN8tJdlr1m9nNpGLqLVQux6Rrztbnm3oxhh8ax3/68S7cDPKa6tz+
0+AVgXIj8EjY9rdbbTMxZyqDKK/IkUBWi7hZHJxuP8Xnmle/NeYkSvDJ88Y2XOJpX5d6F9aiLDhr
YGjz70q+DS4oyAM+fD6rDWXu5ijUwu/yG06vBPm97c/699PQf1vtk9tHkbSFdXE/6+MXR70kR8QM
J+uUUAzY31j5iJkPc8hvn8+QwdsbTEyRQC9AwXzYpm/9Eese7QH3GPHZ3+GGWT+mPSsK5HSOgOL0
PoI1fKYPo+dTS2HatkixY+AxE25nY+HbYUsHgwZyM2pY5SQFovVsDX91gEwl9q+MMbi6tRRsRq6W
/lOTz5ZInANwAEjEZ87ivLC0RwQ6/+9J7x0Fy2kwy8hctIC0XP7Q0rrk0L2hrf6+/MXHB+kRjJqo
M/dTe+Nlw16+Ps/5wBhc9g1r1R4hXtIXtielis7R0x25roadnI1TgHmnCczGwmvVsFH7BFkWoB7T
qmJW6EOChwOM47aB5+1YzXtrAJr/8m3Jj59gIDVpaXoudxhedKcdfo4DcuE5XMqydAnJcD2E+6VL
DVM/rJy0JrB690UINv6QYeD4/dFTSTEhkaCYoXddzGOS+rKojeR991iJUKikrJWjSGnu3N5sPW3j
+x18Rj1cVtsq3OBp2+RIGo6qWEQ5s2yylUsvzHmg1bEzWIOHyIcpawv4tgZ5Rwhc2RkIIhH5CnsJ
QfBUHgxGkTzPO+t1Yd+ZWpTY10hjOY14MPwKSFPyJjv9nw7luAIv+gVcmp3biezAKPX12zbITcDN
KgKUZQrpciq7/gARFhVSuftpj5nw3Q0haKFb0nMHWZLwUxeZUS9DEckT6/GxeXrIikxDLe4iM+Wh
b/CFkxv2a8plUfgsY0frIGcZBEeEgXKooDOwTVOZuq9L3ubn0qKVJXYzHtONJL8k0xQGyQaLZL/L
gvqEyeYCtv9/7+sRzzA7WFnvpYI+/zdmk4dJ7Q8zK/TmtPrplTlicrtWZh+eirL3P2Ay3dkllQ9k
7ZsveSd9vZhZeioKS1itCHJS4UOuYDleS6HrIcWSUI7GXnJqw/wvet8sER1bVwyTOlPNQKpFIbQu
OWhXkLyWZrxioOSD3vfuJTRXd0Z+bhkldc+mptFVIFcjCYno/4xtki6OQV5ZwwQycnJ1x8y76Ocq
XbCBVmtIeRuXeLBItGx3qXiYJHWAfHOcp32fAUeSr+CisFMfgdV0B+WLRDhVZ0d360zNcVViirAm
dM0buGd9sdWGVzCFSFES9b4l5pnVyMf7YEgts8FrLsI968HIx0hCvFbHPuiK8VMt0v+jmD+3xCxB
EmRnqrZDtUxiKnxoW/iVgMDL7+1rvAp26ZWgDdweZZuEbfea0rM8H62C3QnjejcWvsIQcx4CaACT
8fefWm5HK7Uq6vLdEuYJtoJjJZsTfBZvu/5qaufiJHY2hqsYLC1Ft6sDe67b3rKRgmXe+DSFbnvA
oXfN3f9gknBDNT4/S9Hm+OjEN0NObArhQihqq4EgsTLr2eB0aatSgkZHmcJHvZBHcMz17iSey2ka
wRpX2qOADT/IhQyil69JXVOugfYijOBhnwJsr9YyhrEqO58azLyEXtyopnMTbClsTx5Uo1RNN1ri
7RbbpiOJdBdMU35xf44010k4DySDYg1HmZnxQK7gLFkxkRKrgomw55O+UE9IWlsymDokjRp0ARCH
5ilTp2nWRyhx+2ipye/FBmwH0BAhJhY2vrnJmxMeSw21WrZGCCoGocE7P8AWn9pensd1mZyBjHU2
+hxYUwiXW/ATQGcOWzU6s8OdojbFsEXFSKaIwzCUqIcXdk8NTvI+VIOtKn4zxzenTfriPn5aHBQh
2frUTMJTIVZDO1tD3N8JcIat26Fs+DGm0kdCV8pvHOt9TOghJ+D4SqPBEUCBTYBpA1ydBnHgthRV
rxv5E6WBMvlbR/cge7KIOLhut5ZuCnPqQ+ILHklqXHtxCj7RYfhaxIpW/oWDs9X0ElQYxZSo2iuv
kZ/bA/SgJdasB30C9IehZ0xViABTyGskKmIFWlEmbPoF18GRAQ73bBh9cEByurZu2JnyOrMhluNi
JoA6XsVq3l3TaS+XAmih/Sf32QpHINUxzZZMNiCDMcgJzG2icKWxbNY4oYzQKOJsx74yAhzOM7zU
QXgmGvfyQ+nDLlwCwchNpSb42YBk2CwQ2Pzw0AiIwYut3SzArRUOIoOTVZ4eUq49rVv8SHqGz6pR
FrdFtFbYGoWDXHDqnP09w6GBAmqzpvSi/jI02LJs9uHopfcmp4+FGXje6pPLsinYFOE01sujOD17
Wkv0X/HfpMGPY6FFLDKxAswHw6MdnsL0JibYEanJ5LDZOjN0OrqvNy+It0eiKCNkrYtRcfR0hJ5m
ZHzd/VESd6a2pxSUvHx9c8oTcXoWmIiFYwQy7iJeWAhSjSIAdHiyc1D55k9wHk4Mp/CQhM40NUve
H8CsaGvWDqMltF3PNzMGkqn/uTC8BJtio6f8cTqvfE6CWov7z1Eh7t9YzzNeFr2g6kO7l5o8V0dB
/SNzJ1BC3aUK31JtnV68ATWl4oE7Bca5YvNhYiQlVz62GphAy+Q2pc8NV2fDbiYqzqRXs2cfyYM2
CNC+DGa/Of2CJynVzb+G0qGWJ3ON0uS5xUPWQhXvAjKaqaag0LbiCrYYdaKg3ALymbn9WoYRkgUF
tEbX1Q4ENVIMxwy7PRaS5bDKQJN1ATJxWvayw99qOmDgD9hQ9FUTOJCvU1DlPOd3ZCaMwssv5srP
FL1eM8yNRdmynwN2nfd2OSW/SjobibV/VkUP6pXkL2SUAHp1HZn+dkiShWoX0elLha+JF5U5g1JV
4M9z+adlPikY2Eke7FToHHB4DjGuBucPlyP9+fd6vgWpWHp/gh1/OeHKzi46fWxCDtbT6TTWTl3X
I5KmgOV21lYcusgTaTSH9UCaPvkgKRJ5yV0+TPeNBZCgyVtvfP0ajEq5gl3/2uWpEyr2tOPJZDx2
dXd4PWOFuPWhMs7HSXpFBHhwOWDcBZHW8bNtqxw6epV5eMbzvqvrIxr8wZ4tfvo3YlFtP077FA0r
rNtzNQn5MNHAuuITXdjGgO8zZF47irdZk1Xz0600gPYsFsSLtd5haDJ9KKtYz9xt/LGuJikRpSrf
AtdA7HzSx3Rr9tYwFjAJoPr1qPL1yP+JJxVuBYs3G+wwTQmt2Aa+FaeC3lwevHnRa6MFdbIEyNGQ
n6eJwbX+5q4ZSKfCbUsE9jNRN5ejhvMcYs8hoOK1rwbMRJMgjzdzg93TcWIT1aAOyPRXz4hTavKl
Y46pkHNt0B0UilNMfrM4mTjEGkqorDxvYETkDmtG4ASh14yfg0GQRmC3p4In98o/1+qOvdnmeQG5
3zXewF5feIiIuuM9fryT27Tl2SMwZdkamXS3deeT7HAXq5IafSuMVq6b8JbeQUYhVcrl+4dpHNCl
oOMdq+ZZtrTs2yqFCg4u/Ck1JDZyXnzrO39h4PCn4ePh7kFdoaFRCh7rjigIVqJNJrU31Kudi7X0
vP905gUlx//SeYZWK8iXYbpqSxaGw74PIsUT0McAXYdijrK8P8QjD7Wwxopzkqe9wMgvnR0kgzjt
N/vjSg9hOtUKE1ZVCxJ3z56ldLzwkzmLStnC+M3/BLLZrV2Vc8f7tQkhErU+CeBpSgPZuqwiBQnm
rBr7VzSOmFH2UBc1ekujMyAOIxLu4vxUJz0yoHpPQUeFiT4kZrpujjw7XFT/7B05Xhkha3O/tWNr
a5ZhWw69F5X5U0hc8TZ6llG0alBeAJSbOa07u6Pz/MCKoopPX3vrASjzDdwgcy6xn2L0Bk5YnMch
GgJJWv4LeemTK9RuUQkUkIJEKj8HBSJ0rvRm8k6UIgb5u1YTMdwHaRR5tKPFn73XCRszgqvpcvt2
6xLwFg2EVP24AgiX0x1/5H+CRvO9XSUlDmol4jHNcdrGjc3rUeQz+ehsi7UOCTz6UUht6v3vSOb9
poFbaHmIcw/cb2ycepqDsFllNchMlf9AeDjd1jzdx/YIamNgY/HPeMMB2wWUlscVcHONMXJKmIPN
4p7lwgWBC3aq8AeyVdezuUaUgl/hmaVNGhmVzr5XOhWrj+JzNy9eZr6s+QGL3bpHInLMZz/YvAbA
NKPsX8Fwy2BiVZfZHA/ndilsTKtQFBvvFJDhjmJGrQB4GVtjhsK3KLKdkLrvVzaOW/x6QSwyjnEJ
0I/xWSQZRt9Ivqf1SPbTw9JxtWTm1NRkmHukSqiBdgvvfEfqrqF941kbwdP2VnHKjFnsHWB0v+Zb
U2Gtj2xfgx7bz6iXgHjIV7+wJUT/YM1Muopy9SYYN9nIRpi2oqJbtFlsTknxNdesJkiV96t5CoC6
5vnv3WSD9gjDE0i6JJ4l7y+14hPojFyEhwCgk5TkjN+1mnshnUVWEvNtLeheChJ0xsHlGy+jxNTa
BMRiQyqPAMFSzyXbgrG9AepATzbMFGL+jlnyyfA+Hj2PoRQlrfdFlb7rO0aqFAVr/7xsj/1/zOGE
gWiPoOFcsR5EFEaayWlJvgKE/CsirsRR4DsKHnf2B1t0FfzZaK1krEqNvbMPlLaGXJoOowKxVx7W
2MNhpgLEjHV+WFf8dqItFyE9tQwGACqLwNivOp0z0i0v5CZEk1LpuPv4A2qQGhJTEmJr5Ho93/bP
DTXuO0leFxXFb7HMfFB5k/nW2xFAmVpDNp2GuTVLZC+8RuR1lbcXCiCePIsMFTu2rcD4bu/OzeaB
d1UWZiQeKJKwJqbGHXef/gzBGUcDDLVpvb2sFSh+jb7/dKsgh7Lv1Cffto5woYRhVt21SgmkAQLL
k8G1iOZkJ+40qxAuwRaJEK+SZzL6RuhyEnOOo1dwOjg53Py+/j0A5Kzsxi/YN27zxyesTOIT72i9
0WNDwj3tQwEG6A4oVUGwb1UwAgsVhcPd7b8lu4P9Dz89G642ClF/At70ujd6tNvsVx/YehgTjTXY
ocDPp/WtJoPi8tHo8xV+noL2pDhSfi0BcFsyc4bJnU1YK60/gJgwsrWMZ8tsKlC7rDZSRYSPTg2r
riq/u4QjkimMc3gx1zr1igdLokiPsvgRBMwk/aW9JVx+FBS0xIUqz2W8lT32ScCkbZuUNxpHc+Lw
W2aW+7VrSwHUN6OtRBTSHQKISk/aFTMgGgDVZ0ZZCeNuxCAyumAv72Y/M8JLtGzWPfA6F/wkPfZA
KeayajstAbq9zumFz0FCGp7AtqUYFFHcqGlVhye/U2k+uRouQFEb5u3SRtQMmGiROe2hGXZlXQv+
N7QdFr4JHzY57i0nbwoNDSLrl0QoNkc9HNUKwFl6TP2Q7rDHCLLy7DYi3E4kl3opopHfDSM3WSJ4
nkU/1e6A0XmV4x6n9JRFv360t7CKWW54Y0N4ktby0t/6o8Glw2Dyq6GmYNJTezyRSkIUMwnIS4Ac
W5nZESOUY2Vgmrg8ygX+uawV5II9FruHTFXz3gtEMyg4PIw5mU2F3iSyp4ogzj4/Uxh4Ju963RaH
zy+M4n7nZvq6SS5W+Zk7YOfv0eShFrGrMeB0cR4ct8p4/igdOCCB52EtFd5er/aOHMx1RXnnD2M8
44nPMDdxpHj8YXw0ILyiSQOqkfD8f7M0rEuLYvlWRaA01MkMPKCriAwlWrfB1lOwfvcAoFvQzv0B
CJpLLwAQ0Xac0WyKzIYmvxxVSH2NQhUdfH2akRA2ACzlMxRs6Yy9cIF9oDKBL+0m/hGdeFlNFlJp
PHlFmR+cNIgiArAIzi0VcabdFKDFFsVkRehpbNGG+pN4VEjsCUFiM8rnlUuooBMcR2IRCpglvDFV
M1ZHyikF6g7OTNXXNgkcQqJGQxHK5CM2ZyOHk07/Zqu0o7YQeTluk9lz1EJs2nRSg5oydyQQiL5c
aB2WtMwXkqHQxeOtgn+FG9Ce5wP3+23vcES8niEzQeVcGNsOJK/1qS9S9fETqQbqX/8xh/haIB4u
9l/ayKQQ1t5jWKbCPE+QaRo4q6v8pzPbF0q7zn/0EZcXWIBPMbQQ1mz1EBtc76RNMB5ctV80jeSR
sgEHk2pEtho6tZnt5I5bImyM9mYG4um7KGGoKEKbeGFiUUK5/FCF0cjDMJQ8lGiyFj5Q7EgMMo5z
i/cHMZozrQ5EYfJ5fmtAe64/T6AD6NbWvVMq6bB+Ld7cCzkp7/1lgeD81RErO4kDy2U+5r4jQ5Dt
1r1ZAT7ZPxC5Dzrm5BVLnt+VCmGCfx6QncJtTBpjFQ8VpZXqecCaGS+rhVLG71LzJ7aOalaNHLfh
4HVxwVI8H9ztJCaqjfe/LSF3z+3FnimplfYVxNo+PDa1/wdhRFTWbNWZPkh9vQ8PvrYRY6v2BmuT
1sgi/tTasjgx9gkMudeBITbfSN7o+107SRQpxDl5yoehgOf+rkEou210nCkbCBjBBP+yH+BsFsSW
PZgpfHcx5Pj1zIv42Mfx+22n8qAo6UgK5J7TNPPIi/zwGeFaOSVPcoIFyAvjhzGnBEWnjWL5y/zJ
qL8EzDObTMddbw7zlhCuu3eaY53FgAapJNLqobsui/WY3gToyHD+8e6c06aV8Oo4Uf2k2TVysqVp
j19FXeIK+2v8W/ULcETImS+1vUWFrvOLvU02cS50SEUVKORcsR0GbhOCkl6G1uow22gT2G3VLOvL
x14I7GrOLyJlVkXV8IwUg3GdoWti99rCeB1Uu3zRGn0d/XnickQnl8p0jBGw0a8XrfsEht0oByrs
PQB84wqKW8/OsLOiHkadJzEePr+im1NRGyz5VHiJFtztJRNQ04afoaNJGrIvazSQdKy9mdG1qRST
K1XNPdl5KMQgZt0mhbogE6q/rb0+nlXeS5p0gkKumJtOWnrSR9hAeHbPntn7/N3tu35WLx5w8NZM
R4zaW752hqZp28urhQI2AgTY7GfWSYawu1k2UVqK6KWvWYx5Orysgw5lNbgSVwiQhaZD/+WVNO+S
G2aMSvWDAWbfKSjlIh8T6skVo89vcDLjcecXlzc02kKV36ea/8u4fGuiOqOPzcrEULRnqaXi4qJJ
g8OMVlOJnOmBRrw5r5U0HbIwLqlI7UBkW3UA5yEb7fmxlXlhOyZ9dB5mueb5gpTIzUGiKAhqzuRK
acEjbOFTkZLEKEkC5JzFr6ODkqyLCfD7/yoO7tBSMMkBjWOAUGfSp4RfJEQu+AE3SLSPfWMmdLBl
1jr3sodFLQV1bvp3/o1nZ6QEqUdNJUpwbwpb4z7XcR2IDeJ0PADYOq3yhMVIynQc8+bimbSb+c+L
wdz2lfzi4npSgH1XE8CpbJzKtKp/lojWmDyrHNkWreV8WABnsbC/FuL/X6mxFqqY8cFbLCu3A1NW
azPtVCssco4LX5BiD6wrgwxMIumsC4IZnEshPK3a9vYvvMd8MR7F9Weu7R+lGqB6AjHVp3gt8sjH
KeBrTHSRgg4+t7AnZ3AU36r4sQOtuLlPygVG9bPK7ujpnG2j79neHdMw8eBwqZcFKh+KtbbrcKsh
jTiXb5RQHW8T+BTH6R/D08r2hfWnzm23Qafg91NDXj7y1/ivp8PkQx1pR1A7n+cJOlcH0VfpFTda
Tm5SeHT95q9SmfQpb0eIv5nX0JLr2ZDOO1uHDrQ/xB4uvwpcL4DqYVUEbMDBLF+Zz9BeXV7zRgeQ
mZeiVLRIr8cnDuljTEGumpH0iIUsJU0Ujdv4FdcOM9uSCBVKmrkQRV1f9BSTMCWJLqriGmeDkBNH
2STr2pQakIJcrKa9yqxIq6xLantNpXPIC76GJyUHUJjLCWLNlIDc9WZi4WQa/Yddk4SMMvigVv7J
qnPdmXWJ+qnomARaipRzXP3/6fFEgJi14DqX23MJo8ad5uhjyxy0a4ir4/Cnlu4CHu/nWoUyFlXE
j93W5ouEzUqxgJsCnR+IOwxiLIZPq34A8aLWpBgoBmNqtJ7NRjotCDUsuUFqMMNTE60NozCcKioq
CMgpG2XVJ9HRjrPP/J0bJpN9GKC+LKstPd1xE3012yUTTlECBlqgNPrOyBC2TG2vKjIg0+Zfvkzs
hQsdHXWsVIMnP12YbNgkzD5Nv912uEuoby01hhsakz2GXkNic4ws6Gsjl5ldVvcKuRqDa89lfweg
RirD1Jq8xx0iJ/YLcT7BJEn2HhmS/39fvSElKZ8CqXan8ajmoc74zMe4OyoHdpB6O664+S8kK7IZ
GkAkeZkyb3lCxPk0nfZZaDdaEBVvbb0D0ud9MPbUGs+IkqMyl9Pq5pHUD04BE6s1iL6FKB8SPx86
QXH43o+KVCKwa/bDa6g99+60plRyCZt6Q0763SD2yjpAGneAFL2hjPjlu265NwXdsWIe3VXW/rnn
BHoM98SmKAmq4Hoq0BfyK2nzzorkrPJ3y8IQFD9nffzjYbq+xJap5mvSk4CEcTiH7v0C+yerpWnJ
vez/7p6GALqAxSJ0LscjEenvhJ/VPh/QM6xWd1RranqrRnKYi/gwwnJiwJ58Z9uxRspJMFBVXMg4
gyOK+5iG+vJJ3pIhgYenioiyB5zXm9KXL8Z5ha8uaJ1I3Ho/ELz+i4C01uTmbNK3fu9augdo+1ny
5bg9OmlrC5uIq5qQU4MmG6pmFgmMor4Y3E3ueOzNB8WeacdX6UNCNLm0++cKLE+MyGBoN7NKhQSA
lVuV5C82tAIsA4mcpx+9LKnrQekS3QPjAJMJ6ZLrNL6kZWwzejBBcyEEUbY1YEGD4TOK+xfb+TJT
tItmsaFnTzMACkFb8+S5+kj7JlU0g+C1gkfItEtsoSl8HeUslt1altR71ESuf3VZbCDNFAFknvbQ
XXyUQam6gWGdV/SMjwPK/Nm2eowFi+9pwy8jKh35ymJmoJJgn3vfh9cXMxVMhLdQRnx58P0sos2U
M4R2CuYnrhdrUIAeHlz9jbrQcsGydwo8H4rM1Tqrp5EzToIwyd1OfV2QodwCuEFdjqGy88upSUAR
8bihwjA3bZolCHQ99OZwKgRSi4w5WR6XX5udsjLPEKT/fTfz0fKbsukocnXEXaaOOvM+hkiRCcXV
4dOwbTFeXzRQFv9++6fz2V3YjFGu+UA1bxSjKp1OTotd0rmipbmyc02yps9An/2sCsAHGZly/Mvi
Zer7E41Cy40n9U9j7+hWmrpSZcpTUX55PFgZ81HWQIECgvZF7gJRAmVWd1bvKXUOmWtLGUhXZYG7
YaT4vBh66zmAbFFPYJbN5tXcpUyoZC2ImMeAeICFdgupfQp//mmjpJSX0HITvSacgTxiPUXoxQv2
JNtjNk0Cdb7HQW+DKFi5QVwxyDK1pfTnVQB+ieH+mK7BCYi6E9YM0/9PFWY/SkF9J1Os0lVYqFc9
GEqAmmK3mG5YTHjcap8Cmcx88mQ1jloOSqtlz3JNuW/zbuXqCGkag0bx7AvlFCIMf09eRhmsKMQG
iZzxs27DgQoUl/CDWoaIV7dfsKuXgQH9/StbEOclzHtoGx99n56JLVDusa4wATyKE6+W6ikQIfdc
/2rz0HOZ6AzNsJY03tbph5w8fq+m+ceoL3aTjt6uKhiMuUwkIuS4zmYZSzqLo6oisTRralGhDGBK
LKrIvOekQcfXt26TgMcqpN92cZK7CHcG/shYTzeVx4/PPKOp49zITXdnITF8/q/ICZl4l54QJxEk
AIDkL/9GyjVw0Q/dEofqQK0WOSorv9EDUf+1MSFB2O/g15iKvWslkClUpX99JygrhMLD4or+J2lJ
CpWj1XS1EzOsaIANRq1RLBYj/HepJYX8VCNWpGDIdrlZ0kHVwmQbNM5LWG6anhMAK5iwdashwp4c
oaxc45poWzCs06fGeqBj7QVsWrHAcEu4JgmsuSEdipvo7qYBHFg/QP/No60+0Br/b4Wte8uWZkCU
FbNpVyvPxKPlF3Q/kF8NstaKqPmtkx//pZKYKJAYW909PaoKaCuH3UZlEoXkwjZ3vYDnnRn6upLC
7P3m7EmptYj+MU/dkcrh1CjcUFhANm7pec/A6xD6AJ2ua3fsMi0JEkaHCqnOi/VkAQOkbe1W2de2
TSfr0IxC8TeQiJyEza/EuRGK7b19ioI3ADQMqf9fmZmxWgJUa/MOjBO2Ip9M57x6bg9GGKRVL97J
7Wv5TP5k0xHn5+Q9Ym0xP/WqM4yA8ee+JXhsFNErJhzWGH2CS3tEjTnyWrXzykXJ+fCAl9DFsPQV
k61hhNv4q+hFQJctIYjdLYZnZtJY2Suk+n+qalmqEBEBi/K9OmIda9uWjEXV99j1BmXABLsaT4sj
PrTSkgCJhq/JY4yIk4T3TsrmCe4hFSEDHe+xPb2bXkWC+3NGW9Px64Z+oRRtpTEclXXa+0WtIA+Y
yelgZ+7hquOogC3qQe3T+ElR1LxsVur05gJz88A3BJH2mq5pNtgXGTCmys7HN9mZoRpEsA1iloxX
U8qnPhbVy2K0Zrszd+HIHVu+EJV3+rCfV2VFjIOlKsgqOiQoJXmnD5mjlwKNrJxG73qeezKtX59O
uZkJ7Prf1E5jl8iwGeMEYQ2I1+16pmiJ76Q4+qUlC3bqRJ+ooCGnWImPobiO62kIRSIXoc5gMiMo
TySSvuWCckuzIs1FgmBMJOkIsz25lk1fn0PyHKYljOkABQ0yFIQ43OEctYn539LlDQMR9TLOCufP
+QYTz5drOyXX5Yd9IgDZX6GCTDfXemySBBIH9YtnfewmkpwrjjlMZncXqrYXdk+TC+TyB/BXC5l6
ncmP7vbG0kNWCXDzcvR9q9QVk4eWIV490ZgJtEzAgsZ5FAYPerSG7MQ6DzYtmYJxeK8oWYKFe4Zl
JrLt0GD3k/p4CDPKk9Gg7A4UO3Al9NzUzs8DH8sSLEh+3YR2wGNjSnDCx/DU64/l+GvAFzo2Vt8b
M+/7sL1yeFT4wKTa9eT1nD6GLplR4QPIn0rUKnbaQVmutnM6yVaiyWHE5Iicwk27hqvCsYKhfZdW
pM4N8qCUpHBjq5DX562YjkMVFJOrtK55boUIWHCWN0QRY4nG66w07dkbzE13LUsXRjrRsGtjYToP
c5cyEtBwv6PzznYQWDFWdsp0c6WlYmw8I/CbObATkTT3k3q1wzSB69n1sbcUaxZJBsQso9VrIwL2
kft2KBHMl6XFFU3Vm8cA6qDT20afBvtTGjgfA4pWrjtXO/iUI9zM0cIeMlrjWY9v33rbx1Dv5xfL
EOlCOR8AodYE3KrTIFbyo96Q9avs7vvyKZxCN8YAtMDbXTeIGPLOaceUmXYIyppvkl3qFrxCRR5R
XEnlZnewqU9jIEHTz8GedJ45QmSEBViUUWJjqyZDMYWKgsynY5rlHeVvK/veGHHS4+8idqoYCfxM
QI0ynNlUMQff6LIlo/eWx7PO8TG8axpPaBMbPckXbA4po60f1hCIF/SX4Ef1sX9Zmp1TJeI10tcX
7vTppu3iHLdvY3ZPfPNPCWJCM5YegngqWSASqgUyb+YXJQV/vGoV2W8Avlvb8zzihwwuTE/f16BG
3L0PWFtue7zi4yoU7EyuUrLIuMXFqXmPx+IAuGwpPIrNzciWfO8nx5NZ9FqIB7j0F+W4qHGIeGw7
SM0q+24zyLGi2pOEzQq00F/QPWAvdPVa65zJQGf/GJLQHEvtI5/3NzH0u5KUpfXqVja9vdTa6YWg
71Fn/WzoIrTeWrUuKzK7AVuIxSNe4wG3wO8OMHIjvjW8Et4E0xK1CeA0sHgaXudk7ELT9uiGqBfQ
hThT5hmvkdpU8ryYQSsDwR1sOB+SLbHy+oXwJ/1UKJ+kl3XSOiwu6dOx0Dxxr+MZdkb5ePUlWbZ4
j84AIIb5m9OH4GIz0cuVVPTtlIYVM1LQL4RixBgYiU03xlG8dFMAiek4/ktgFlfE7LeNORrxIpAF
8515gFTH+E9p5ZQ4WNks2GTueWFF00xtOrZNN+sDpEqQkaZfmqOTmhY2+2yAfZGetQbJD6g5VolA
iS5GtPW4ZSy2cDsaaF88rKb9hGNVglnI23L70h/lu03DS1vZXH4alXg6CdLpUvQZd83w7LCa0uV2
NKn+2GJ+MOWANd1SpDJ7dNo6LAKstwVSAeGyVF8bsKSk0ywvz3AYtF7crr5JaGjb1QPjlgoiDxqi
EIpDI86I8c463ZRvLIVgmdXGtirFkFNnNqVxjYmixNKnTpuviDizzQ5L4FH8hOgocRzxD+YomKRz
5AKeGSnKBjdSmY67TCPhZz6zmpZ4ii5dWGTcSYowciS4fdCLnqaQLhCz8Y2J5ci0FYWPSxImz363
jUoBAoC991C6cDVIlzAJQTwiMtHav2Mh26SXO8QT2Num/Zy1eV1GQy8TD+91sTNosELlBR7aAyxO
uidWrUcYfMz37mmHZRHjDmarsjefb200n8zC2ieVAfBtW8ZgmsXYadwDTLg4G0gyBubjpFwIELaW
9f588O4Gk6ILjNIFLCjxy5l3Uf0+yvMQIMjWsc341GTSJ/cbNSsGt9e/N+LHER7XZO+aKUiC0t0Z
RVTEjMm4LvcMSJFyEbPw73UDgpm4Dneaun5D6VkRr3w+IOUn/Qjhwe7prvJZFiEzyOubDrLBKg9A
CevNsIlTv1Xw+TGGeo6kYnszYLf7+FuObafAhQeZk29EpM+Hae3bKLXjjNlwKw+bKfRAfvg7uzPx
xR3o3A2JBccSRha+KPGFNc+tGUJp9LrteQmQb+Xr8QbKApPqD4XDVqEggYPdSAj3thoKcsKyXlJz
XDaJZDAi3VYR6MLOp+XtqeDiD/ionyzpcRC6/H+jnOnMS2+dejMp19Ao0W3UVmxrX2CXT5oCfFfs
wb3Mq/kBPnouIs4TvkRtggaXUHygi0OlVeoTubFCxP5gN0CQtrweMTLdETNlo+wi66ry/UhYBX0j
ldeHu1E3G0hn9QkXCFgzW0xNU2Bw1VoPWnuv59541a+XXKkDIFHaFcHmKSXrgV8VDKyU4s7LhI0U
YaK/nNGWLRlwf29O2xq+73uXjEToFJ61PbIgWrQ1T2+OzCy6lACTZZlytl+K6rYL7HT7EReUpQPH
GEpLnXPOGZYH3ocLLeMkl94MxZjw/jjOt9QcASbenwzJjUppedS+vs3udVTRh78sGzRcNRqQlea3
TaLHzeguVTAnmcam+UkdVo1zPxsebRT4ukUpME8FgG/RBdXqMogC8LS0M4PC2Z8dGv7Jnd8VfANx
RDK9fAqmi1A0OuPvKAzxAQ+xhNYxr4KqZcRcFxmdb+vVwFsclsyXghIH9lZo8iBJDR3eNgco28bV
D9inqb9IKaYXb0P4CSbjVJ4sY3GGxk2UyPLF3hBSyENH80jcFNbNChsN1biSCB0zYcT15IdToB/P
T1XdIIkEWyVbYMv9FCf3Ge2u+3CwoJdC3y91YvXhjNwMJnYmXpCLF47gRyQHA3eszCXHuEXfg3p0
IQlcME2vy7lBwD1kqkqz6OjvGybWEIz7wvcAAGwLEjs5Wwcm3cTVdoCrbZ1MmldnldfUbGwVTzwX
ep8sF6WJ9axtqmDqkqIb2UtNSWUWATDxYpPz/EF7yMoNQzye4DS6WhKBYezQxjHwFsagz6af2oum
RKmAfY1L91JNwpfr0VjVsk/xncHpakQ7wt+rWaQH5sVu3rgDHOUyil5G63hdsrOgC5sHfEjSr83D
KbVLQuElYacGwciQDjUUVSzPfOf7O6ZwE9gAZ6Ht6Rznlx8/GuxJH+YaHaO6bRr5O4zyWPGlhxX+
zQncW9m65NIFXnnDbe4iKVI2ZcIF8LUJx2Sq6oepoJ+IYv9eEEnXl9XzrinzHgjCCymGptUiH8TL
a78HK/QcgNJoo/1VVRJrgp9ASBdgQqULvUv+ECPQpbSonjsQCW0xksLnV4cMRixU7+zCfJA1s6Fp
pjzf990nf4UO4UHLLkYYtgX8wfCxzzu81pCPP+ITQXAFEUJIu0vXOh93W939E2LaMhUaQJk1eOpT
m/8yiYfOtDzdw45yV+TN81CUj2R8ePk1i+2fiaS4JYHvYRj4lSYBCLKfl6vCJNeCA9mqMJUA/6Gj
YBXfeR0gS8Z3TJxfmqO9t60UGEK5le0XV9zOY2+RFQjrpRHuS1yqrl4DEM0bRLgCAb6w2VKE+aoQ
eoEdZEZaHg/n/6u7RXpAdgqZ8tkZkPOkmcBYQgeFDqrmykN3noOhOLY4ehaLOxLRw8z8O3LYC87W
+4r0P4wTOT4Wi6XqWt/ysynFSVd9kOacOtaRP/q+bg1r/yri9ajixtMxcMLCMS79Jad4D3Ogz0k4
oG6LF4r8zpZNAU/YbjLkUu93paMghuwOnT+zjif3sOc0oKNLDz3Uh70a54631uj3lbhi26NqjSEr
sJ09Annb9iZtl8MoLMn07rvpR3Ke5O5hwTIjhpm/NOIN2+LpFUp9kbHAa7x2oaCoECDT3IFqM+h0
hL8DOYadfGHq6GmtZiSACLJOrte7MLiP3IXF8UiCrxnPsuLYc7ZMiaHywBf2H20FeDFEyP8wzYKN
wBl8XgTjF2LUe9LhcwcRmpoVucW4+VbZc3zPIp97lTcbCQiID411S8p4D06QI9XLRP/cF5NMMdiB
JtB60Zb5q7spPnRm77Nx6qBYbq8TegeEaqqM4ByRayup9nKixXmV6xZIAHI9gUFy7l3eVW4wcGVA
8cx+91hwT1W5qVzYLK5Dwo/xjtNpM0T/tb4fVLXVnjOuV/9GEPy8eXcX1ToxzZjdy9CzIeOOpTfC
LE83Ao9q+hJF/NCBui85lNiLLTOSXhG8Yu6zfEWkwEUcR06sJ3X1cN78t/+R+6mzOEGsWUvZD1oI
AmrFb06lMP+hAqTCzw7pip7YAKfy/3aobL3qTw2aD9x8hzxMByTVLA45J4NzBPu+j9owtG4n1G8s
b/OOjnLj9XWGKmCbpA4/GaqCvKqMa5K11F4+DBS4/uvx2dd4nVXn2jh07QaevbKg6BqtvgE6EoPv
t8eq169bjrz/2923RIYxfdy8zzfPpE/YSZ/dC0FD++80hzljTzGiYyC4syd16sJRWYxksU92d6Id
6wuFdUf2+/POd4ooeIJLjGrweYzw3YN8M0z/H1bE4nXZStJXJ6UW2tzdSF8n7Z6Z8GYE3IeubkkI
g+qnaccDb+DsF72WaG+xg9O2DLuMUtZoAGfaXWqGqSWCDTHRDAYy0T0gU9TqPAKCQPnkYT8hbew+
LlQKOM9tJPOoXYqeeWgVMMl/pgm3N1pzSBSzwc++aBAnZxDMryXUJ5yPwb/wwdDFt0KR6ayt2vGV
7/vzuIMQsw/m7YbN0ga2fI8xggGvOH0o2azofy9lm3/rMyY1HG67xLp6qJPOgNbj4wJnXCsPMdKW
isk/WpeHhMf6ejKq/TmCiEecdwE43T+h9vvcEpp2XZsyBVhzXfuqP6kzo/H1fiMevZ3n2gdvxlnX
lZW+wtQAnspoGyO2DqHi7sadGs3imWlLkZf3GccT38sM8tW1nazArGLrGFaV4b446QOEoBimhMCs
R/UOApNsjpDt0nwtlM/uzef/1KlG6ojGkfvbim/a1pAuLw8djsGYcjyQimL8bywhhF8EmQWDLfRK
Q+ANRNxtA+vVJpjQiTGthtR2h2PzXUUWlpoMeURXx+a8ZsD0tkOrBcKakS9SFxe0QO3qb9MoQWBj
Y5T0DU7d19ZfkKI9tH2EIjyuzWAtcMFowK/e9aF4IzlpRmoc/TmuxusCy7zj5FH/KLm9ak4oEpC6
7iDeTw7I2UD78IRsugRgAFUAtA5xCi9JfGx4dEJmcFN6JAPw/Hix5Ir90bhSULbpXckWtCXaBCKx
RZ+Nm6d9xnP4PsnWb347DUVb+swIIpRKPqTUvrrlouCsDmaL7Jj5u+xtLiKiiMG+SF4CO3ot0URc
Wbq+Dr7QNsmw0sPZoe75FcjmFSuXcbhM0/Ri7jn+zTrY8M3O4p7clPa6RoJ+2GR0D8ca68nvohK4
FQuNnLCRoQ5ci/aRK0p6H5cFHvSYqnuUFUmJ4Ppb8aqr8uhPb0ANpYDOua/pBRTy3mpuEJd98jqY
XK/1ZfPvaEujEtqg6hDC8YG8uXDl83iSoWdhqRS8RyJ1jMlYDrwHc8ZPynr+dY4YO+Etm7tSNZEs
BggdRg5aivaMBSxSGD+3GRxFd6XSlJDuyP/9tCcygZ1Qe9bTE+S/Tpx6LaHqdeNehPiF4hDHMTiG
aAe+U8wxODdkK9g2JPhpJGVFoC7I9cdyq3cXZxwuYGiJwPtkQqzvLI3umaWnU8rygeHRtNOi6mjV
sp44fQXqz6aZQDB5iaLtJ81F6cVF3lun9ES57YYnzulOvnoWCRLm8vL48DjxCVHYQWWVP3orGRqO
kdZrqRoFEtSfEQOZxeQkYIF+eXQaQCX8DILZ31XfhRfiRFUe1fERDUkbgVLSvtPyTPi52Ta3Wu49
722ftEYNJ7GUFY7ZcyVlo+53dQkBnzEQiSBKVlo2jjv2jc3OHPx9ma0FlKi6TFog8guFEAExf4W2
mNJX3VAfmUCMrrWhio96XsX0SdHDxEKFpC9m9viz0od1K8YrbX6/9uWsr72yFzfibUpGWv4iyEiy
NSSDjYHWe/3q8+zK6MaodxIB3+W7vKGORScOlHkHeU26oRsGiV648PmIHq/bitqVCBDs4xI5wcL0
GgFYzREQpIcXMVvLQmtDLV1X8jtUXYQsf3sKJVDljaiFaaTJlaSh3u4uVQ9pr8n8gRxAp+rjG8RK
gxvaU7mvbj7N8vaM6u7Vgr/PEDoMLAsq5de+exeJcTTHHx1FK3GCKdTRcnctwnyzZm9bE3Od8XUb
a6a4HSS+f9OJV7o3m9hxpygA96C8KIxyuM4EJIV+SOqOKRRyYi+nngdZ4tyvyTarrmEHmymPU8Fj
rGTIysycsHHoAlABpy+ehPIYVYmFRHtwhhfXPGvWBS/v5QlQ1DMdFesTdZe9B4lROnkgd338w+DN
YSpoqdcUpUiXfJB7BG4+pqCHbYvR2XZ99Kb8I5heVSMAKZ1XTUbUhzYfXVdkGlFlCV14he4mpiWP
mp3vQs9rJsKXeRRh8ZOt6u7EaF60NU7G3lboFegLuF25iX2qjoAQcxM3Vs2JB2HtNq3ebKrNZFFg
4g++rhyexsxgfvChqJQS92d9NgvR66tpKZBewwLkWYlVQYgLEXH+cdeZIWjGgMnXwqOOOYX/10nK
Zc5/nv8j+UlcVoMboIjeP6XhsJuLIOmTAPJrXpDmbDEhXdA9fLTMSDTJAYD0yFWJXQl/WdFJL6Ud
rjuA3hQGZM9jYjy3tt2d6t7vAIq5HQdt+cbwA9skd84N5uigeW5S9iBhCa4p5hWuLQNTtGVXHMjL
Pn+y/pVNKmxu5DirJFt+EEFUUnuCXQNa6TYWTBFjnmJ1vJ6jr81NnT4QL6f6zrJLXDJRrDAEX1AA
+9JbvFtWrPrAgzOFQZNbmTTrNorjBo1U2e0sHGyqYUAckfij2j8S9CMqcIhHo0YbJjHGNrXdGaDD
+n81AQVmFSzJhwkiCQxx6V+Ip3mn/b97lzWnUbGFIMayQDxceC36UQx6SxekW9wJKr60iD2GVkqS
42j62qQERwi/MrpzR3sx/FgEYzhVpyIXvpYVK4T7CzYFWvX0zOUSDZ2LjqIcsyL1RWFsCz+DrDlg
T1AjdjC3zGiT1OodME0RSk5MYc/8fkJFRQdqeCYLSkgnERuFJ+HMv9PdZCGKFb2BwHKqExGOlmGc
uSzM3AyEqZ+MWXPDlfW3MCVu9uXEhQPGRsNG1ishsm58e6SXjSJLoVDXdvcOXLINv1hs/8mP9tOL
oudBcI4BmEtcaW4qe8sNLdIfk81TCN5NirnVOCdYM03UgeFHkGRoD3Tk180AMZtC9i8fWGmPbh7s
eKZzmJ9FeCci9oZ4RTlmsB2iNAv3HUtNQQDp612zN89T8mRTI0F/G2X7cv6RJ++dFeR770l7rftA
+Gfp4yA3JFH2gHQWgrCijjilaWgQUXMumCWeBw08kI0LAHvAOg/q+JNv/2Yx/3NaY09qqIxCyQSp
dZySKPZVSQZCuPC7ySNDhWE/i7RFhOCO8/4wLxPrsW6O4uzmIQ0ltVvSw6izrt03R+9Fmx6josMx
P8ZiEGMSzF4tAcNkpRWGLUM+FNbqvnrv5iQDnCP6OYZhi2RvyABFy4bx7oG0n06nfVIMU7037/9F
wDX4EevB8OP5zZiOfKQ62i2cUpTyfX8SbFqMzEmp8EKw+Wr56namTAXLa4lQglatmOhfx1/iw3BK
iSmvmVXhj4n5oWqRxXzauIPv/UB9HyMPBblTH12Qzggj+T8AZNX5Vgg1KrPwbPB8fsxEtz4wlmrM
RgqTi4javoPyh8Vk1hGD3nTbqQppYrhL62Th1LHWpSJeM/Cv9UvrfwpUF9RVzRwyeTTw4MdilJPp
F1DrA5Mq6ta4p1SBBZ+BCEJkUURVssjGfuApxjho4To5LeuHjKfYjDHXYU9ewwet1dZSDF4Q8znH
i2nboKbw5P6Ke920VPpu1Z1tB1GAyU9W3wv4I0UicbW7k8jWWTKkq+0Eg+slNr6UNvCPho+5TnZb
RVUE5hB5aOn8xSnSZRJ0P/ck42sZ+bmADOH/6ricM2W0N4oLaS/Turh0oX3umaDNWnjMF8gW8NyN
fQvdOhTAuYqU8Z6uKHtDqvb9qDKD/c+P2WkV0awiUOICX5SugmdWZmVPsPAy83Is6d9fQMnbeWSB
cbxXXewTssYkfD06bsN/Tdc1Rtbf70wJiBB+C1HnJSMmsOcMjoNI7ebZ9NqWbHefh6NdrCiK9ev5
aONPKWjIlJ+uaerJO7MqRX+S2D3BgKPjMbT+1BdNfj3XBA7xGamYV0SRbg91fcvQjRPIYxDR0kwJ
NyINVrPckaykgDBuS67BZAl+aTsRJ9RdNe/Pdu7huxkQy4qH3dHgVak4l+K+EASjvlzEbmF+KEDM
Fs0STkBfJfJ0r09iLHJCvb3/WK97xIMksgkjrFuP/9UObiix4V7x5q/JOMAUKigq8KUykwJUwHwe
2zp6MAWoSBrVv2sz2R73Dg3um166f/AMUa9nrlQNhodlsLeB4cx+00OZczOS/9aOYwQvLn6ZrMFl
AQi3mbROjh2RsQKVkbCCtW3bnzKoCK1kx002Q7fee+Ehj9DNRgcTwRcljRtjkvk9oogYiQD2pSSi
SXSVfAiBF6K3uNQFrRMMqWsv1O5odlZR687XsnqnmUlX/MmJiPYROYXg/A6VwTxexlFaXOvYgxbZ
/pwH/E/4QCNUmpmQwBsW41M+vend990dhqbsGg3mesL+6NipgmTyHkH2VZijY03flM0ZLxrYGOto
utZEhEPt6CfrDujrkA+7SMPvmpNzsCpWGL2drsWW4TQ9gM1iCPd9/BbYFf6mA+HgdQF2f8nAARlp
1XWIRiXknVEiBajchJRFvDBWuWZU3msqOKMG4jabG4Vo6zTJBJtw3luCT1iSwHWHXuQpJAECBdzV
JQBQ0ziW7qMZqtTybK2k482U37Bw3luatKbmVGIDGfLeu95SDFztPdPkHcoBSOxOJUNDws9Ket0U
iL9WkIfmYNYvkLDqJbjAds0ZNLGhog5FfSyWX0uYoQjwrTsB56UG5uuIcFq7/iWscvJ0PWnk9Sol
3JZCBen/UnfrpRjiIiIK8jtJq6TjSSUMDWsRyIsV5EUgx0lVh5dh/ey2fwkgF/qIxhSTknBN+Knt
kBvvDcPrORhiikA7AdexAfJuZCg+1k3MLltPGDM3bi+IYGrGye6OeEO8dkMhKVhICl8J2cbQReup
Jk2XIx082eoOzYHDWJWysBGAoZC2uyJx90dSJ2/z9mHhPzcuzdlpY+StGDd4hbquIOMaMFZzyZkj
zPcjYY1zK/+pADPVILpPVjo2jLmCxWt+K+S/t2d3+CLDhdN+MzMt34PAv+phoxDDNnw/OesVl3xU
9gX5OyoW38o+jU6LNJWiLJYa1qWOhv53cphR3jzOUS4Dl3fY/Aa1hbQx7FSKtKFM9UG1x0ifMIpd
1Y/Ken/MSKd8sazLcwAgLyJ5/DvijuNJ+ypOR1k5FfFCwmIR1TSl6nUuOJkt69jqLccs3/OTP7tn
6hvcMXKHCdaGqTCnYR0CZLb2mr3Csq9dgXqwC8Eu4JLkCgyIUfEZZ9qj4/CaJT/UHW0uZBAN+u1M
arLelaXTffx1xq6fgPhwG2pMrGG2tKbKdfkWVhDZpDhYopb6mO4cZHDEGlKy7CX/+FmzlL+X0HZs
GzgCxQV9EMnqSbdTs28D8GGZai8xHYesQiKKl4ioWnc+RgBaTS2YVToGIQE1Is78WEK4ha1cLJXD
QpSku88a7uFsZyLJ4EudD7YtbcgPWJaSs+NVbsMqu9sgW9+1piIqerElGnAYt1LOHnnQ0u9Mqu3w
rvqJGJmEtrXzwMd8ENcA70spfURr8hmWXkGnmBCRFf6Cl6OByqB5+FJ4jtx3dPt1EUchtk0Z1QLH
qWJLhuAuR5/TLLkqRlUYSg6ZUk/KaJyflbscEOvczc73KPDwxtnr+y/Svrwqy+1MbnL6DAgi/ydz
ZHOxjihOdIJdBNdyY0q7Pl2WiTP01RdiKmGRd3UoUTC1eUp1He1iUqPwVCue/VpFbuI8LimxB+ZJ
krCSoL2F6pneiCd4YaK9J2wYDXPePJD1K+t5ZMqarHolS4qcC/nHfyUSW4Z1Fa8+2SGsaYLiHF/j
F36PnAICM/5bPYPQrsmB9+7FXV7s71vLMdsvTKOLfDQnZjuf9/vo4eOJwakH2n7ys1Touli7oUZx
546vQqJmmxUVLVZ/kEEp45uhNzRJOMffT+C8A5fDWOy6SNukQjdhgzh9j2Df+lceHLKTh3gJlA9v
XxlGwCRwmVOOFkQmFufdcEKK/spnOFJ+Itkh2dJ1oehOnrXPDWTw8GvV7982hSbIoKuhFV6yhWhu
4+rkId01F/FVRk7y00fwd6w7avsaTLNMskeX3y5muPqChfyUee9tvCzqcW16ywqz6Wh9H0vdbHYH
Pz5xiU1oZjrB13PH/9deKaGtF2kiUblz5mHnswOWih+1oe8NPGAYZpqJk9GDgYbGOdgxW/YU65PH
Kw7mDYJ0U+XmsDJsxcT0Fl3AzRl7Lvic+JipnRf8Lr+/vjSZsmCdrvtgA4yl0Qs28esaRIsoREHD
TuYYYHoZpgkLIVjDG7vOh1sVrWF73sAzOQlqEuS5ZTM65aLSMMdS5p0F3ByCX24OpJohj6R0e1Zv
uFXdnDr/HYUf1/f2LaF6OZdlzFNYsLBprdcg1H6plqwed16IJhxLa2OFloX4mKbqTjVkQmX1gM/P
0r07650DF5jby84KXUNH7Kty2XQGp98uCFPWAX2v/eOUWqr+2HXiZhF0cyCOTMiCnN28EEm6cAvv
pAm/6odD2oPbFEq2kz7RZ2anwjx7f2FtMQhAdQXiIEnoGmrlWciEPRaHgI1TCGYeDfjWhFySIIVT
8TB6F9xC3258IV3OGH/V0LDY8MeQYYtVIlIOvZt3jNpxYklhxYggJi5wsZ2sOUGOREDxo9aysRzd
F58FSaA/mux9iJbgVQzlw9LDtUNSxpjbLkaW70sRtDnSzf3i8io4gdA4INZcjG9TGufbXLcOfGPb
vvbh1vRqYUt8HC6KoO6mrfBAOtBE0GCfNejttYYIHiC3kERUA/vBYt1sIJBmpMOoJJx7hTbRldlY
Aqk0UxvtXciTO9GTqiUS7SDYnglCQfQjVOj16csSC9CdZzsAXQn9xy6BU+5gEvc7LCe5ypfRsTBS
Q785nvISjQr60T5rjQ6WJO/79Shum6nsFxVYGEtHs1/YZXwT4T8ZSOfM7E5RsRrf8AMqiderhlYw
rqJR8Efn59qVh7eJJeiTtBx3Z54e/f5R4j4bVrfdbFEVUWeeZ5wXBOy4rwoZGwpWuoL8Gnbx+jyD
YdVGfH5S3J5EHZA1ciz3oDkuqHKELfUYdAjiwjz5/kwpL348TJ9FroR3x5UEmy0CNGruA3DHKzYE
RYM98cY9S034Ji06F8YC7JttzJrMkI4H4DRPjPTXskHWQ92O0Rh5n2KkjiaT9NAR0ThlLwnlF0Vv
aHU4piKhkWGbYNCZMkT22Y56YPJW5q5UGLBk0JFtlE0nOBlLuZI4WWC5hsVk1bSs1efPybEahX+A
0TO3uGFWiwWJOGsndmpado5M2LGGci6wgphXfoM+k7K+om5Vz6QYvH6A8MR+V7ru7pXWwPzhr6wb
RgO31PMOEoYbt1SMvqKJKR1Du63WGGlMOg/NvssC8qj1z7k2l/xw0O8mnMYxaNinuyR64WxDShCM
mqHaES0D1WZhFiMXQV4eron5IeUUrUHdzSsVBZmso0t7wI32bORonVMhp7Y8OcgbcZaJ6lzWPjch
2fOnyQpxfi7pclpaEOZ688PWyIEaiFHqNxD0dD/kxacx5nxT/9cVpnPteCncBVrO3BE6EPK8IJ1k
RpPw5Sv5CNiMk/yvtp7lMXNF9Bp/k2vJpVjR+v+KL1bM6GJoccAotPlqAsR3b7bLxWl9d2Ad4RXc
4+6j1fhZIrW/T7aVyNHD8nPyiCfUUb23IozArJqvTB/bmWW2pJft7Dj4c7f00Q5nYx8gzv7bm/kU
H+p551L9YebyjPULkwNuRVIhnvpy0scPu12yxa4Bqwc89PzIpB1L29LCzj6EedftNgoBFWrCyxSw
dp9SP1sK+14nqGnDZEC5m7tAsdgxqkjvoiCeaVVUO4xw2HEpxchkpKDcH+eXmEtl+XH27GD653mK
Cx0gLyBpJa5ry6fFqHRNjzsOIfqdBu0+STkCdUWqoWz6qXQy+Akue6t0dlex96i3tnnwCRFppL6H
532bAqmWPgQOQzYONkwPXISxQNxLB32lG2QDCcTsUsbu8llku01zWRKjJiQVn3MCB1DF7pi7YYkq
54Vt9jVTtFgQe8TXgr2OrX/RYqMPhwUlszkOuoQxfjGUmSPTeuDDpmc46aK2H3RFriJMTCgf0pfJ
DOJgFbe1d9YN329YwY4G0JUEA2ZnW+uL5cp5MWDUJdZgYk2FFZcCYnHrWXYGQPMoMopof6IER2ww
j1nNKDqsFm8q92gFYHVwCehzXXmDUrBKsnpPB7k7I922rjbo4mYSgmdVboWTPFYSBC2GXcCldUVC
n2eaTdVoU9LGtEN/7rYsgW7iF16cnmydGYGkV7/Q7SB+N9wOmUDoFyE/njaENPOED93z7sAjwjKl
Tc+gyNPdDfWMMvGJRRgHImzL1+Eg/O5N+L7PXF3jzTIfmRnkDPPEh3wGfzrAyMVIuocHAF0taCvv
O9tzw/Ht2+oVy87ZJqFCYHeMQ/i9N/ymDSjuIwjXoNur5riR5DLymBLrSmnZB9R6Xgv6FeluSGvU
bwB2Mp6/GwE+zbl9bMrR/L2y7jUfiI/0Ym1A+XfMKvhODXWQ+w9zpq5slUdMszp7wj7WilK6Iys9
0O7MsVuTeXG99PMGgFwV9fkog++jBEmPwkiD6XMPzKgggC6OhDdoZgLW6Tjl9ALEk7GKSDyDJtRA
V7zURzmwWNuc0lYnexN7UyMZwR7BTzhQScTlk5csTmYzOgqGpZiEOxZMl71z3vzqj/FOO61yrswj
aNDCfTVGrwXU7ZpARm2lC4j5UAcWp3rfogfISfobMPAKtmQppH9IdnO4Ke4m1iPYyK+rlVjX2jCO
3uAB37ZvGKKvzucL+ieH1PDMSQi6Ni1Mi7IUQYimcXXMZlVopRNjzFk4Sub+tjHB/HEmpQEiXLK/
z7IdwTPSSgRoy2HxGTZgXYagx234Gn0io9RRI0RbJ9s/jKA28Fcqu9aKHNHhIfcPn+w1PLF5o33D
AGrKFE0WoXFRRGzCxmqPX0o1mjelQqxR+6KR0UzwgXPFzo+pQBeo9TcWRunuTFhcac80sf+ExamU
7rXcWKgwAE8peIMk2tHuZuJZLAA6cXfFXY9zB8XiDd6SjE3XTyuJvz1zJ15hgcIOEcijiwNfbVRS
jH50u91PLHulHYy5e6Qxq3wt9ezidng0C/CrsXD9bWnMjpEFucJ/plP8oHBNhYt2M98NN4d+Qg4T
15tRn+uj2oGjkaQ/MUvgD6jyeg7kS+9R5hFTidE1H4e0wTXMaSC4PK7ia6+kr/urGzFtZWpo2Gh2
mgnc6XGYE+RGOnchierIN114OH0+bwOFoVk/h0b4isnwqyXq3dDFo2AkrVqi4f23+/7xo3+zdMoo
Y87+kKPgjlKiu0M7nk4S417Aq0xtUg8jRwDEX/S2se4L5pdQAlCOacvOR9u0XIHqjkPLf+bB884c
TqPrjly5nqv2EbqKbaKTIekyz3DayauYHvirBLV72j+3NPHqkhk8FwtoYdVxKMmq79xPjCTpAvMC
koWclsFk7ix5ZA4yghX0snaBhe7uGL2ysxj69azCpzzg5xSfmoQ9c3NpTTVjmcFavxMR3Dz1I1tN
s61Sz1ia+UJJyF8HZ7dNCH501qudVhyiaQ7U6wzddfUGniUt/Lj1KEJSrhOvSGLYJ75clMyB8Zlr
wUQqyWBHJJzxEb+lGK3KGmcMeO3HDiQkmxOAVDzBgc5wNu0ojF8wsTsSLa3k479Zn0A4RTdosjoU
4cJsz4Vjgs9PKHpgiaFJUifldxAcOSwP9mkl8xSUMzHNL7DZKWKPqyc3YqaNM234208nOLrlvXrU
ZFETVhSov9hVbw5x1nmdQULSOyy9INNMx+r0DqHBU8KvuulRfPaCZOIwZz/IT8/3p9rXICC7jKEX
C3+l+YDngqfTINrbevXxPCmGQz8f4YzCKXKSunDiqOHmo/356GDjWl29RHGpL+mZtZ6ydIsicTyo
NtghBMOKgeXbWufTn1+V2gmRkmm7yTz8HNW463UXQQoJlmws1bHK0KrOR4VqWwVXu3h/oC4xaxAT
v8jzmkI2dWbbYYwrX+iW2elLEhfzSQWXPKIcEpvDWOHHTMzi57Kxv3Vr5ivz397T/1iDhOt32+oS
nqszgPbTPfo9iOeLuWMNz8XymIp2c4M4AqFnGo73F/IuFZJmlnZtkBDiPakqhtkXm+7NSkP+r2tq
89C5lBrdHVb6p+BLuC553mrCf0bmc+X8YsxPJptTB6R1XA/Mc8ZgY3lk7IXzZuKdu79OxSnhc1Ub
i5jTEY4BSkwLbVXCElNGFIseS4uHwkWJLxGNZw6UyEgvJJpMPpvHxdqo+H4noFUAUJekoLy8ApE0
zlDCR8TetnzXjlMgoz0K4iW/vjQZ+MBC8/16Zvcxv2FpTJoasE3KACg9HhQYeEbOA2BMb6iVFJ5M
tukLjyJiCeN3KJPCS4LRSXqYmWDlf1VoWnsRotZvUs671sGv87BCG/TF82wSdTzHUP9P1QRYeLMG
b2KTBrOM7utbdh2RluQAwLF4CC7ZgdntThPaXCdgs1H3/6hCeXdgZ4J3lsIzxiCzi2EQ38K6WDu6
7WovMv4GRnMoqnrML+ZtNBW0ySleRsvt3ubf9KD3I//wVVAo1pTWI8mGZPg3D46G2cE68WW34jnK
/aTSccpn8TZYAhPmJHDjSICuf6O+lqXKaoONZIYYA9K2zbhGvo30iovnSC1N8I1NwPufRSTbJNSD
UZpu2B14tdAQiBf3M/wWylKIdm7pcyyVCdWy0zmTxyKb1p9F9APn3O4L9CgTE7aO1fOtHddQnBcQ
XSPmIRZ0K1ybUAIGaa5xFSEM7bPvmqdqk0Z4Q1UnSvWo6GYnjYhoE0LbxYlIiAyKgBKrHPnZ3AEN
0ic7lufs9gs8maW82HCOH0gK4J99q4xye+CuPlFM6IFhrLbn5IG0flmxrmpj7J3e6LOErMcCXi1v
cNSOolguNJRpHpEUwJWLpXeUWSGhCuxz6/2GS8UX/WZcg0sSIUzroMUr4DmIpcx7cUKu/9e3AH5M
zd/mxCPoV2u5oeLhlgcZxrGGFQ+pShv/cYJLzoVoYTKyLUtBrCmznp3zmxOfiNY33wivYaZPxgGp
uS5ve41G+JIMtxIRKpcopc1XhZGQr7ubTY8Ml5/4NLw1It+rGDXEgh1f0pmrJh0OZs7gUcBfV7Ww
pEp2jVmhnp/Fq5bG7jUWwO25m12Gkx6JAOa53PSnHrY7BtiB6y8X8GQYX7tKiGgIY46sB9kslCY1
VgAKt02LjhfnCx7aDrbnQMnm7dTljRCUpFALDK9RsZkoRS2gXLR1CNpL561eQrCQkGlh84h9m2WL
j18UAq26DESZQ5SrQZ1zVHXxAuSUzArWXchJoloTV4oyL2MzqcqkPQaZxqLSUI5ZmFqva3M5QYFF
h0JHnJ6ROWUURlCbqmCO/ZQN21aperKgq/RWMbOwbVyritfT+StPn/bbcfVNLjrdDSsNAK0KrlED
dDMyp+9TZPi5Idd5CrvGnvijfPduJjKtAHnnpcmoxa2sugdmyDGS1E1FXUzsoCPElSF5TeB33CSq
DkiD4ZGMaZ33eUjKfkt3vmzQc/C9oVXU42BlVwXgcgQcf8Qkc7ZP40Aiq7cYLDu5bkIPTPvap7GY
kK1B6J/0j/DZJfxriYG6zNCPd2DidAGGk9jCHCVeJf1dHWWRdpwH8Xybf2RCcgImEiM+7kEu5Fi8
YuM1JhWyIo1mSJaZHxPEoUiXSiOg20uvJsVN9X3Sa3LSm2+abegidGU84FSMVujmf27OlJhJylgv
C/05E5HdEjszGCeoxubWqMW3TAVdAulNzpD+Tg0ghrJaRMBaoxT3sESLQ6lV0N1bFe9tHIbaJUNs
T7KbpE59gt9ZkIux5yGhBbi9ZwgMjawN7EBngr1EzJ7LEpOk7+vw96zRrtxx1KCyy9/VPIB9Zyru
WLEKP+OBQlzkMa5HYoRlL0XoqG71modE+AbrwFiQXRdcBuaARXrG92ZKdKry627Zl+/db2XwTlOU
VienODpsUl2JNcoi1nozh+YuLNCdInQ352IW+dXSCVB3uikO7/NSalNf+OtGFgnDO1ssy9L1PT6u
YbsSV4jYZ60+rcx1+UvOMtzSgMGrhyBahhqk2S0DDGGX2AvYpP/vzsCl/1u9uBlo0jRgYhGKRrdU
WUH+GtYmANBy0dvN9BlO8mM/JMOH+hdDMbyjyCFa7vT08daRWVDR3X1RTd0l/GR+deuAgr3B1/Vs
zQsiCCuUSs47Bt4GXY/2b1CdxXST8+zqUh+GJtNe+QTwekOcmSFJpG8CSc0Tf82UHRW/fOD4VPQ+
MMV9Z4eVQl66lLQACmH9AD/HqoAFI+ezgSZCmQKoecmR0ZiRUApD1ScFHp00fPlNqXAR+7dI+d5A
90py7mlhFMk4+5WyNPiECGCJxKbw5fE/IHm9dOX6GFgs5beHnFoBKi3kg+pR/5flkSBdruO7EdVy
mFZ0PX2rXa9LPCAAnoc/z8bCwHO5EAjzCbu4iUNn+6ukYHZ2yZ/G62eqlrfi9ZpNoJvdST5C4CL1
s70sC+IFzVXjYcXHiI0tEsfwGkCyWZOmRIqLAZKyj1a3TVEF2JZ//n/HAkqv8PXUGONhy0ypENxT
Q5x9pxwP1EJk97PEMPkxpwT0+XsHDbb1y1zOQktGeKPkOIeZygIrbiBxxIQvokK6lHw/8rEwGpnQ
Peh2LE/f0s46eSyPn2XlqgSpO6w35L7juFIrdVQRjCeLb7bS83wpvwRrQ3frfiljTQefaTL596wM
aYKNZJGFiD7bBtwBly/p3PN6uYnlxfrF4BYNlm4bgmLtWOfMqOvZZMv+t97P7CGDGwTL/u+SlJ3F
BD2Gw07Dy5qHZXAku81+41ieU1Dk9AOS9YD5yeUaHK5nLlICd1dfDGu8mkSPgyCY0dAzjV7rELjh
ef5bwOkz/lSsQvJV6LrIlcZ40KSnxrEqPu4ZsgJjlWhCB9Vpgo8g31EJIFpIy+ded4NoiDP77XGZ
wGV9pjMTFLY28eLEtMHCbKv6EIE6/z5VzacRhKXOcH32/70gySLYMklxUf52Dbk62unF2IXue4Ej
kfnWBZ//LGuBtbGfmTtndVxxypBas3Aa769gA4IzjcooSQCkGCYY2sErLdi9+5oYnS/hsCRqfLJ/
BMbn6xIaKpsAJLvTb4WJt4bChSahpXxKsXixBsRH0KcbZvBYbJCSjVJSMKa8lqpDQ1yBEjJWaxRh
uHTlfwomqyz3tm8JapxCITqPDKG0irqxL9S+oLoWjEfKtCdOutjvT3jpXbp8EuKYBEMWZtRSLRK8
EOYNWc02/RCRI4vdv8MmZ1TBTwSAKsQ1P2t/5DIGzm2nfOJ49tyrugRfbJLzWhHO/pLF4YjtInS/
k1YhRtYmhT0wXArIzO6qN0t8Yq5t//GRVFFX6w+6TO70y+XzctcWZbUwf2agWcS/+z7oOE85Y5qe
rMaf4uTr4+8SRP8JFDvTC+ZP3GZOLi3dC3VMIB6mirrutvhW6zShQLbni2qxdlbhXZmx9x+xHG8q
pqrM9REO8szuXPMqSWVj76Gk9gOyJlnbZLHASU+iIloH+AGA9aEkFBxjV3ms+Ou/lOt6uIk6nGh+
Rvfc4VoHtA3wcZwEAqm4gxz6lDF++QpxnFfkjbk9Dc06oSxbURuw8u4MFl3kulEe6hk44HU4C1le
dxM8ofuvstzF5fmGSAdSfJzfMvKTbjjslK8tEXrGSPB7zROfTc3ARHURVNrVDPAXH0gXtqtsU+08
IFnvj0kMnDraTPyM6xqMPmvoxqDzhZE4+kY9qgCM9822Jt2rMIJFLldOdBTH0H86UeGAq3Pge4oh
RokpnQoaent7euv3qwn3JKPpLPpIayeTwGXLIS479iYT6c8NZ5B81Ui9eI0yWth4MJFV0k0yDS0z
uF4fhx2pMZ++V9HUNHBlKkxgFn+p/k/xKuVcNySh865c82oQhD9RhNpjOGyfS6XHUJPj3+CVirXg
V49SP/PcU13/B6EG/+MqLRSPmE/4+WdcPihvJJ/sLQdAICIG61GcWyCjiWO9FEXQbuizJ7ax8Jv+
aT2rbVj6hIEla92qSDetxQGHY63iotwHaU1ju9vQH7zTUJD0jfG+iq86EvAC4enXrLbaSVb+6eVY
KPMXvQHcJFnf5500MWZHm29v3Fp9ruPXA3W060O1H+N5KbgYWivdaq0CBJwsifTnz8LAEaQLeRNX
4o2ryWh/MBBi3lEBLSzNn2h5H/B7KooWbgKcoAOeiBNaejJ0jKP/WOcTH7aCbav26XOlxFAgYX2s
dNYMMeth/INjJNvo/+Jdrnw/CrcdKBNEUoiYEGhWGYwEy4SioSfkc1aEpSNlZex803gcNrB5f04Z
5LprjGJRYoUzjHC7D1QGNlzf5rpzx7LJjOEioF6aaKPLi2Lg/E4ZRXBYgRjP7VVk/c3zYzDdaWcG
UbYTwgVAVlPDW5hRitNyhb1WFmLOqjEdLSWg/cMIcJO+tBmJTqOZv5zMqEPxzQnwK6XXmRb9b8wp
4MwZM1uubb5dqPDe/57xbq2jaTyuWyfvwICN1mwv1js951xujUtZH3X7scTo/pQfO9hAZzjBTMGz
+ADCF5/gfwnlTPFwVkoKg9lOEBvZiP+F/pvBnPknu5IYQo/4QQI567LQHNePypLKQvQarl3D9kwr
/npwkyrZcJra4B51VWMwyZR47BX3b6Q0X7TAUWutJyIgEWn5K8RBxfvWsQ/U1x/XXIzcrt8ad8nW
XqGUCuJkxWZQHMtj+2g8mp0ptLRTG5yu/Y6T0hvvysEzBhUZWiJ2thSt16QuS+sWMLQgi2oTR077
/7lhlUNQ6YcrlMIH2CB3eB14Xob37PONgosbqpJstVs7SfX3G9BWNFWXhEdxXi/62VeHF2XANIkL
zuG+WzLd+sBwtPa65l8H5FtAZYo9RxfRdEPQ7Vfr8BFSkGjgC0cSVrg2wzbzzlxGZkcP/S5I0LwL
mg8dwgzdDu9hyeQFIXwo+H79fSxlkvVbKv/bxyFmE0NwsRnzwgFvogwyj7eXI5TbsLnA43dN9uOV
jTA+mJXh5zaMD/V6SUY73b+NM4IxzTTZR0+WXbjuw/E71f4RqVAILnG3pLfSWQD+5kZlhiWUCPcR
d+EIbiOZN8P1kwVuZDezt80fHFnGdboPknhJ3TnTtO1154vkN/tkssptKF05ZVn7owudXizQparp
7ho48f9NqwV/lJfgxq6tM4CUKdXo/k6e+um7M7XkZuMVh8i8zxYH33KyNWWiN2xIr1t/osLZZ8IB
ys1wnCOtfgaOYvXROfkBdu915BA2wbQrVzVF9KA3NzrozLQvIllCBj39eUYg+Xc/GZ5HYkBkjDzW
0fGv0X0iHVcZNyz/helYiVwMB1zCA38Bqtze1/74nh9W6XacxGaZgxiL8YRo0zQskUdP0tlrVN/0
CXpLtonAHLBWwf7nVM5p/0kyD4iuFjTF+C/ZhwUffriedlZf94CMBlP2O4CYNvoKqy3hZInZJjZr
9IdjerM3Ix64l3BS2GmLOUT4va6298VYLAxLvM2Wb/ZmDfbTWbEMgTFZ5FM54ZJpGlIKYbZ7hwXT
hx0GOt5e832hDQmHhaAjg5C1cGFq73ILKP5E7Gr+8dEP14yMc7MgciLVeIFNHm0RbiiFwpdiIdHz
F04nVi0v8AmGfzs7tAFwqWdVTwtduMA+epnlEzROdzj4BGGwpTjNx2w8ZVK2gGuNQkxoDB7KYG2P
aZiI6Zbun3QNy4xS4oYtFWsVv8jO9X7rm4CSt34NZgbO8jl5DgFQJrD6HQf756+KvKPCxD3WND+M
tHUu1X92wAWnV2ToGZsnxNdZHlwdRmH4QDELPQ1RutTmz9gGMocn6318EPMKumiGCyN+5Lhy4TCu
WLuG4kQzVOGnoyWZfIYt+ggS6/3MSOacAc0MOnm50pvb4ntvSfav6Z7muoDZrGBplS+vz7tcAXLM
5Cz01hVNC7eQmH/KAevdn5wZnkEeyM2aOOLphAXibr9wxsn9O+h+RA64JVHSYSxa4ujB7GOQrSky
3lgmYwmPtnfyw4w1qvnC0Vd2isAmjyRjWI4SMsIDNUIIWPMyEGHoCl69PKRgMTiNjG08W+aDVTra
sM5WcIRSXMqz6qlF2HiS+QeBzFiCwnFOMk++YHDUnIdpAGS8fJwbsa878M/B0JanRz/uz+biIUDy
xCUfP7lvnfIX12AC7dlInfMddEkM8VH1lMyg4RKG5kGsywykJwQOTLkr2vsP/bOMkQi2UfHX2nsR
4zmne6O3Fly1cfcKexH/jH5ojyfQeXhMDXFGPagCu2cu9Pf/5YTzWmHfW+1hc4BICuBCMU3Y5Iki
dUHTTE6PrO50fSWzc3t25pU4YowADwZQgh3C7IyMCK7dnTbfEgRxhVq11TdumTopJ1tuUTZTmn8v
CzloqTgKYEzlckQ6xweHNgQicxKjRdpFi0A9YFITgzIN7vDDzobnx0lBPHVRcErdUkaDJL+G/x8K
asH2RdWfkGr57gf4WblVoxLScGSZ7BtclWKJLQ40xJLzpVk0U/S9K1D0Wf85GKX+mjG0lvNNvA3o
RnARVchpsLPMgmzXyhSJ6HTlQ5Ca4OuscP5CDNgdcGlc1wpN81ASfh8CgxfhX80K/yemLtWaSfNW
IrBJzNwg9XiN0R4giXarjpr2fo84n/N2FbV4md0SnRzKf7hgMRTu3Fm8N+dIaWDEW/8bBC4hIRDg
/Rnje9evtLnSrx/Fjz+yL62OdOoXA5l2ZBcwv0mgWJOaTF1DsoZL5hnMEcT/gwAefMg56d6LmxjX
7wroGgEWEAC9FQkziQiVwRT7p2V+ZGGSPhGBsEl03Uz/ShorkkpqddIL6mydxzCnE2z+oJYG4cBk
7yW9y6K7sSoGLLhC2L5cxqB+aBik3xbfmTLDvl/YZm6A9c6jstTDWpdIoAtJzeFsbK+c6NE6Ct81
2wAQP0KJnV5AUyt+mRnBq593jgvYH0dk4Yfx2cXFyQzznQh8HCK1MJOt3qaZzVr5AyXaMX8gkjwa
oUaVW2MC/nzJ8tgzp9rPuPItgBt1rryFDRWw7s2IJpxKYW42blMRqTJLnbll6sFm+H1j/lQZW0Vi
rrYCWB5uVYqLVcQblNCLI0NXuw/sfdEvIDdBrzMMvt7kLmUnaDCSzdemP19Rb2O9j3gh+601CwmA
ByB+D0OoOCufOWK9D4/V7StVzgr9DsAcij7A8egkDBtnB7N73uBoghu1vqeVcuYzkOikRx+DKnKX
Tu1IJ15IWw2ECJIhGvymkc0+dKu7CA07iKiwz39Rub65azM+R5J8a3og9dcqhyv9hM9CMYU31iAn
P/ukhkAo6ogVt7OYvyK8+Uv96Li96SPBFD41upuTdBmADWLxeV/fuHM/itna4uFo0BNvrJOo5abu
VMVN7+qdP4Bl+BFa2nZ0HPoCvtAJsTYrqB6ElBBjXBmdejiR/qaZi1jqBwUcz/ITqq8fwk37gori
zB1CHSlCjy7H27dfRuZ1FRT0cL3zPPNzC5SNTtFdO5fSz951FKS5QhPsvVAG3i+/6C+ZVy1X2DNA
q8UoVtBqct771CdBOcO9XX2O/kFCECA/A71HmKN/46pTdFEEsCu1dfyqgBL1jdbwAcArYrbki0gT
uzSPMmACxuIyqlZU60nE+9D8CES/cvMKsLfQdKAbmD4yyZ4YYvoSpYHTtLZiZdJ+ejV3niyYZnJa
30v+9uVP/ASyE5f2XdsybSuNXUTDMgKaUcJFp7c/AgfiPId0pelPQbuYO4djUfGSMu1rBWU448fU
PBRXd+AqbT/wf1Wc+6V5fujt2x+WG1Oz6FIraz945uWFk26u/6+LNTtrGv/zdDNYt8UaP6d281WG
RR9TqSoaNtZybQbtyvxb6YFjTan98xYjqIDYYkFX9NBvdZ11O4CLX/eTgh3snRa6fiu6PP8+YzS7
BsjL4r9MJFfqyUFQKhA1AUi/ZWyEGMSkCNWf+jEC78C4mh6pVh2z2ZzBp3e+ROxEKDVODA7Klx5B
+oa5mIrgMdfdgtiJ8PKvAWuzmDjN8rNYb3bjQQZaj4NvPp6YzSliFkhJiPkQp5xio97NHg4BO+u3
rt+hUltJpV94OQ7WLKkom4ABzLQ//7+/RLBvhzwZiS4a8RZRm5yHrt+4qP+VeBxJ3FoCqD2KLSyu
Xl59QyjrlWPWncvbLrszJQ5moeTDDQiyK31KWha4e1n3/sPxgdmg4rJz91jK1U5dimBOmW2FcNu4
czugw5Wcnds5U2p/1YS4JD9guOakYwk4WD900JKLrbiY4GkLFgea2cfRWL4sQlv9RNf3PJlQm+Jb
jQxSnZLFfXZEsaTntpjuGPAPJhtudWQSdyP1x99MsL/JIWcFp+wjseO3HFRwvq2uP8b3C+k0QOQS
nAUMZtjR1h3KZIF5h1wzV/8SSlusjUR8CcB9VAdb++rPNOCwY9hmSYDNEvj0Zi3QmsBHz48hCrxY
v/GF+v7Fi0I/gtIXeSlTS5ACtt6DUFKBY53zyfnR8revLUvV3G1VLd6EDUCA5FCOopCmKdYkxWy2
WyI27kGbrIT+DG4aWCf/ZOo+0oczAOZIhDSqZSEZywSSHPyczb8MhylQRLmwY3vuN2F21a8k3C16
U3AjESLS/BSzDinQEvzT3qOil4Kom5po2FJidQB7T0UzNYx9AxuNbwd7jbo9I+MF5qwEASMu1Ehp
EjiPwFZyQ1hJmmtHcfUVXJBsOssLxaK1mEQkMKXWzxoqYoPD1ax1w1SEIgYJtwZcG/59mKbLYMQd
M4XfOxshXNe651bJOvne6o2PPswIaASMNffcXWnP9GqRa+3FHoT82xJiwnZVd7Hxlycrv1QFkqHE
3cmuH9P0ugBeeYNiK7ZAk4rmgxDsHV5Du7sPKwUD9+jX0cir/XbddUpkQ8QJXzZe7CRfgt4/Cvsg
TcgIqi1c3GXQx79dnhViN0M158xzpDHkAbksmIu5LY4Iy/gy8xQ0rqdIFbxZnpUWl0cOrFL+uP3S
YfdlEyOtVClUWWMRtJL2w3JiUHkUZodYgh6ooYQWWwdL3mySJIDh/Dx2lF7Fvif2skzSKW0RUy8+
FSPyFjLE7DSnCAFujRzRiKKdtZOrRIJ32qN2G9ljJsc0pe/UUeARU0UHWpreVXhOxD5QyuhpAxHx
ADkSJuNVMSncQvbynqNEL3OS8axVCZCo3G5JPxQOX9UAqy4NLWbYrbIxdyEIYIA0oqengo0j2e8H
c6h5HIgzsfUi6GcZI4ZBRBuWNBVc65Y0ExPvqUOofJUGHXmr348wZS0XL1ChiNhc9PlVKtC24wnV
mLIFCcomhzzSWPwBGZTdLBNZCGcWWwybKRjZqkfnSe0ErWRfMSCsARGuz552liLHkAQY4yvvSyMv
We9NXa8KEcPazo4tcnIL5j5q2ScQPZJ+eKSXTTQIjwTynpqmNKGu9cgNMpB2Ql2suN2hA3T36V1q
UTPdDrq6/uz3ukJnXhNx0VNuZD+SqeOWXDfdcwZ7JV0lzMUfNx70eg6q2z/Q3uBmCXX0u57u2fn2
bRKGGyY6FFlGybW71BX7Uh0xN3j6myGJxVU67ZAbWLJB2SRSwS+d33GLllfVWM0nrNCeBufxrifk
VHxzuehawBD4QXYDoTnhA0ZYq//Fgc7cMLui+IqLFBRLfZzcAkg6p7pEvI2t0di5SHragoVzW04a
Pdvl/ZX3can1lTlpHSP7Hhv47wfxDAshED6rPByKr5/kAI745DlQbz7+0RbCGeeIIuEAHCZnNWL4
IBOnCUVpkKwpsoZamSUJn1mXpVSZ8oJwqpbxaAKM1abw51LOO4+WrfnX9xS0KxunUCFZpFLveti1
z3ayze5UI9vGYM1KLkRnBIGw3JH4+ZNb+bDdiMQd78xozIkk1GaWAAB/BmNak1b4qtzERCGQQddn
qBRCOiYTRmLbnZVVTX5ns8xIZPa8sWAh//VCEINK75T+FWuUNUZUPbQ06m33k1rVP4k6xZVoullU
2MHJAATJEl1wb+KelAuWFwqKy0MJAiIe0NvhTzqIof1puWgvKO4fKDcMzkbfnUPSUxc9JtCT1s/E
yYx9Ts/DdN/HqM5q+G9wsrU9OJI/qDLDgObSmPTl+DNV3c8MOWReGDVg0JslhRUoxEJJnajbT8Xp
DbJxlbCpz4awW7dUvH0ipEsWoxyjr4/ynkHhZS72ustPInvOlBshOzJY7mFm6TEXqpPESmiJEKDo
zrMmiOeirTTz4CQzFA06M+xRpfKimHCFyW6riB049VM/D6gpdlS6orE9AFqKiExOlXH4Bv35dAq2
O9dk1xomQf286s2kNv6emYOTPHYH8P9+F3KozL3eWDjYfFH558j9LqP2uhPFzHSzMWR+iLB5WZci
Z7fW/UEVMrSJvRiyJnT28fRzwRzpdSTe2S/MNzlQtpv7GAXCnXxkl6I3ZJu1OtVPCDCoJUaPSWkf
D1m62znBRAQrKLA5wIbOmyKMpQgaUBofVP7jn4SSnZy/YfqCgiIba+BIMhs4zNLro2KkXFletqAt
LOpqOHLenYBw/QH9/Y6z998LQM4nIjfiQ/E86VnDMXqRZNUzE7goh+XWrDXZ8iD7t01X10J08cvE
f27/TXfs6qqaCiHLUq/9Unfa/KDZzjIXBU0vUhrNaxQ1cmQtMN66GyBoCq4lwFcFEzncyqV0F3BU
Uf74fRe3UjKoojj7nGSo2jBGDoqXmryeJP5URC7IYmLowEDioLAdC9Vs+acaIOaUSg5HbDVVJLB8
WbBRYonjgDcAFqSR1dhwpI4LY96keItZOMTKSYVqu+jgLa9iJMT8/UUyGhCs9vCC+G03gVt3oFmt
KBTBw3rzGOJFPzRybhMU4o3G+pH3SkhXJJFbJafO29OMB/VlOP2vZWYXRf7U83WWILH5ZuLbO6Rj
PlthMGla3FcuwtbxcMf9hcDgYwlIxi4a8nQXQp5VuY9KIIzY7N7xNjYu4fVlm+yjYsY628xs1W67
zp2Ra/EQcr0/WOD8Ykh6h4yWA7lsL3yeCK572BXoYja84hu09Lsp1TnRnMLLElMAo5Mb8yLFY4v0
7iBtkzIguQXL93K0zRyvQF9OP8bDBWY3WUwRVYMWxXTfQSNaokrjjwu6sfpgGSAAjNJoDxQ3ZetA
4EgPqOsHyzetqEPBe9HqPmybcA7u7dHiblUSxLOo4k73sexvdEu1HY69oGgDqIAfPptGVYaB0Ix8
w9LVSq2BvV9FXW25W6oKcZT3I/gviDYvN1DNhJuXLKTSRpy0R11HP4Si4dJnnQjLHQKzT3qvrnrU
4iPcIw4jIyIQiqfBqHCGoQYyNjCzV6/xiQx9QfNZlgcAwXHpG0n8KZCcpfxeEpAhrdDnezA49Tgx
UEv0HfHR8orsBc4GkD7BtOkXvokhVtWeffVPKS5ZkKxJH0U3xh/OS0H/3oKV13ZcE9Xg9599R5Uq
zGwfkGrgtBKCQqKb+U6ggsQVgVmf9u8wleHlGfzlhNlpX+4rDmTazuclxOUlWSyrT687TwrsPHtq
QnC3yIrCZy/VIY9TH+AWzStZ0zHXtD9oDp9jTsOHN5dWymlv6cSJGvuClZvQJGpc1h1HPzl9pRCn
g/kXZMn77KSmsEgyBUqQ7th6c7A4zeYNSgcVO+0+oItJNOyDyrW8SbOiDXCnXcZRclkWSgKCc9OE
7Z3XKiNwdZDW/jDUWZcutUdanlDMijblmTXRWnrIsJQNg39sAczUbkVS1J8LRqMspp3tOrVGm0us
NuDfsL008Bul2ibzMg9IFiryYsj67UoNwUK778CFqzlZ/L7Bbyc/D999b8Va0RYmhN/srt8ySmN8
NVlifzV7lVS+1U3TU0Qecg17LJDtKQ5M2AzMOL4km2tLjdZffRf1pUBdKanB58fe/7iH4BUl5m0O
FdzG6hWrBEKk98xuwpiN802tsn2hFuispHRjpXYrhC5vWvu6Z8tjD/Ur8/EHXCQOUIw46t6rCzWW
g05PniJty1pouIl6+h55yE9BK+6DNKHDAVKOmAAKQWab3L46z7DGi2jGvp0Ocp/A9RZwL1mt5m3u
n22UFU8sJlmmFaTRsNbh0ZiWVFJvFp8ogWWsF68pRRjrldGHZYsnvRhVjmI6FT8Oaed8VtuJ1qkb
5We503c7FLTaYhUCRDE/XJ9hd6lD2f/2yNzSd41dJtyQiox7e/0hRkGo+MNvQSoEeCz/xi2P2KMK
Dl1b2yMzl11VPcc7qu7SUJ0kdFLnROAzdKQF5J+14D0veo9YrFSnPyQjGZKk4GrdzUzAf4uPl/VY
cY47Rjw2vw+GtN8nu7QF4cG9h2wtvRulgJxmOWE8JCgoXZlCqrER/usY12ZDlHD2JRWghSlrLjhG
qwfL048HGtNEyqRJfOLB/7uQ5lV25LupPqZfYDRuzw8E8PFwB0nLZl3Yh3US+eOq+3BswP2jiyMc
XuvrwcSOq66lBoQZIIyYxLbArNEmjx3/hjcidGjAiSgvWacfRXnfgYZNvkrUoPmyk1Qf4E9UpRYq
nZNC5dPfRkp10b+IZYRjeEAjRcx4RHe12zZtvI+43RNpkt6dnpzqsnUbnL4diitA9TeljDe/bR5B
mMMukxEjVmoGAoW1jmiwaDgV0oHq3XF2rwsfalCU8Pl/dNbAVrYFOq9v6FowyCk1jWHvd68udf7H
+vcGLwt2FJVn9GDHODutBA3gX+JSf7DmDQUspUmA6oaVRi+bLfAcPNczcwU8CbBXBrpKCEy+Hh/f
e7mAd6rjEuNtHRafdeo96QosTKMLpc0MrKvdSi/m5WW+sxSO3sFyWXWkDHTHZz2TwP2JRVtODfrV
g3CMoGqeZIEE4Nm88MtTgHNXBAIRGYyMhD37T8PkVILHL+gXpfom3hVVOB/6MRJ1AVkYn8FTgqZR
lTMYHILqNL8CwDX4aIhfbcQNYWh6/NIsS6BseXs4Z7n4O5fQsXuvaoih85BIQendcpBrz+QSVaoN
cTvGCjbF8CSPmKJ1F/kO6Qp260YYHOiqdCUTr5NxQ7nAj5LsVUXo/7MtPKbXv0DQm4MTR+1va/O0
RAShYuC8o8Bq3Dn15XoePkGdijVwARi0crQs1G/6Qgh9ltjklXJslgCFmhdtGXfRDGLRgabrrGGE
RO4JGaom2m0C2KenWTNV3u7pAnOqMH03eh9OT2/HIfxucea/ALnDCNXudCLY6YO4RwJ0H3cGcvf1
oW4GjUOsd7q7lOYr0SBoZggxTzOAIJqQ0R7hED/o/sfXXnSOQDBwluZtyhkcgsXPwwCVIrED4Gc+
wqPhZNB7t4nVZ/4wFY/mUdSmZJZhm4T4sv+OCpln2/GkZyGqlsZqq1EyD6MN+1KGcLa5wL5qI/3x
oKdxTwrJg3FJYm1wHRdMO/y2rs6Md/8C1Oncwk3VvJBt/5mUW0VERPXIkraGNSEMKScx7CgxNIkt
rYfLd4v58WPDGD78ULmwsUQfKmBjDMHdC3ja+AFCBu4snA2ngT4kb2pd47pVXoU/uADpV9bqx4ia
oJv8Rj274A/0KwXMvydFLP7M8zZGXlwsolPGrjZPfOeaF8V8fFYfNVMyOGWLqENQCYp8Dkgq/v/b
9/Bdte7Vm3/YhYpkp8XkOVvR8b6dOTqlR6LfH4d5wW0s/dSz8o9iw5RyPTRh5/YTyrhQbXEpG0fv
VIH5DV69KQjlup7g6NrH/BzdxHCbpW2/Ehav3VuWqAaF5ZwYW6QMGF2J2esmlqX5xQjChK/Dv8te
hrC2t7fYlSuKG5uvqDgPF+/R1QgO8L3css8PPBmRy5pNZojFCr0mAVIQnE27Ya+a+mW05erwFlAX
SQxR16aCw/diRVeSTJh8ogypG7DxtuQcAUAJhMynpRyMY16gTyvVhEgUGQnR10gEAXtULZkQ9l99
s601FutXMDL3ekul9XzCqcrmuS3Qmk9E6Vp5CppHFNtu5qOdYNn0KN1gm81N5zIZeIfwZ8Y23Z/2
4aZoEK7+WDvgGFwNDpFEZ0aiP0ezlp5XJMojUecNKOk0DWOfE0zTnk44+OHRoW7dkAdVJ28ENAot
3nYhbnr68xggpgSQUozATZPomVz4bJAHZJqLj1s9wkpV61RIO8PVIklAQ0kcqPZt+4bPBABmRz0I
mVjqwRngVLOcoTmIrr2PsbalHhRBghJHrG+iF+jEIHKK3rblm57TJi5as14COiK7L4FzPI41/bxE
7Zs2WMx7iFlM+MV8u4gHM+SaJXx6gICwUWlojiakcqczzbzhqjikwgD5NuguhYEFW2sd02y/+zGG
DQXNaCzPcoQxoP2t6I92ssaFEIx8bqaHtGp9mWfDdlPwvS0uFhkkjskEqzQQ4+sl82W4I8zxJR+V
ic+ygxgMcYuOnXTwTAJlOGzoItHdeWnYgMPJvSZMrBKYKoIBxnh2TGwHMGz8UDnJ7sEV/BJL4M7d
Wjd4LYJu0FSzCjA6zCpEzIJzwrkb+p08BkgRnL8HRTU6wrC/F8s12Hg19wP0CuJ4r2ncaWNXaSDe
9ocwrlTy1BOVTiy7sxda2VM0yj1CigN698KiP2i5wXZCGVafKL1gsuz3E3cii7aRPinhE+6ErrvO
iGWqKpITzb1/2j0l5s45zxu+TjoZ5FtT49MQX7VE8Thn23BIuS2u8YU5ABlS5REG+amoBhimOZok
nVc5jdGeXaqsfB+0V7kUTrubQx9H7n2PTwqeSLs7V1K7vIRZNrK4+fiHTWlGHN6GsDu0nd64bjzJ
qEu3dTg8dxj6hBts0DypFYvG1nGgDTgzTM9gEMKs2pRvT/4nGvIYJTrmpGQc6/M8+Z0DTlJz/Szt
ma06vQ2NxIENPHb2ZfRRrsjk8ILVVQqsQK943hzhsEYcTXzUsM08lsZlJOKYn7vw+agHyjy8SSbI
IZ1tnesG25tBEyO52xMXMIRpPW5nHHv/p48IXMu4LxNXPK/4BQmJ9Qd5CgFV/hY48n0LZ7PM/aQO
Zc96jTyCy/fORNayOCp8mS8Fi9voFtFtNzin/Clz12/Ad8DCiMUUyNa34lo1fm11lNzxXwiN0p/s
upa6f3vfPKZi21MNhN0UNFaFfeNs5dLmIn1wdSQmSTsOBDa5uyNVNwUDzfHP+UDg2HmEf9kvvqr4
RUpBKc26BIdRdJBy7EExg6MhWiiKKSZ2K5+eIFqS2Xvs7DuF5Utkl8ll8bzbfD19gcpTLXtmuZOE
OZrs6Op2mznFbd6ukNZIaGs7MsW17i7mjrqaxYFXKrHBJSYauGQYbIgJow5ZQhEd2wWj7eRspF0o
9L3+jOBiJ+KBfRBbVdq+r4/fiY2zakJn4g6/hlfXvXZ1tLkuYYTi+RfGGZdmaJtqXLBF8+ZtRAm/
A29Bbg2QdKR5Z3JCpoxvl59MTXEptbcDnzdvObM5TKRclwBvUAIGJkkJIjzOmv5fPHv9PifmJrNj
a4l18aDJNvDpKuXEbo4B8hjok4B3ihTRPBV6OB0bgbg0bvKkpCtQVbh2J+34BCbxyVSHK0CkjK0I
/sWAsbopOQJ63X7F6O61NkWuAXbby9aYe2IKc/wAfk2qFFPgoNtVc6kaga/kmUMlMKIQCwpDL0Ea
XP46CcOXjyofNMe4ONZDqXPupNg2dRC7qhDD2H6SNJK7odQfNKhp70glJOyC+beaknaj1chSAglg
OojgXupzG3A4N40x4Ag+D7XzNBS5u1PUnn69yReAQDnqsSB6oTG4Gak5ocuiIaAXNbcrU1qL06eL
Rw5ghgvFpyH6BVhjOcgaPGnjSPbV56cwfm82+5q4lVMsLnXn/9kqtU1/Ag9BBw/anaVzVxXTockZ
wf+2dzwg0HRTR1SO7GQ4Kmp1FhHpF3l9xCUkbMCE4/7OUNzpAoZQ1ERDGvAgHCvmfliUNH1lA90H
+u0w/FvTR/WR188ciZ22s7273loV59SrMi4ZNez5WZrzs5hz9Md+FG/9XSubqfNGNh3au55tzT2z
sE8jUsmQy8jJ+qULv3cDGoc2haGQ6Mb6gx9jIGJg3hMIEviSglmawaO2oWWkM2Of8IDxXE3Ndpro
JrMdalM1Bf9POOL4fBtgLA2KbLLjLeJRswiGSI/gTGI/SKi0y2eLdVcyESzYYeowlC93f2z+SJXk
dJa+2vSAbgjfgC/m55Svzi7q1xpROVETh7ku+5ILPkNl5b166Ixa3vm5avQ6+DUzpfuCWmfzepuA
1+aPQ3iSI+gzD9GAsXgLZIaxnRC1nt9YGXrZzKVVam74Bvjhm3UlG+UIxc/Jo5r0VOLDWykDlNPB
NU21tNL1InQ4PN9Av5xoUNyoc0UTQIy6Egf4zRO0wa6A7CUjgXwNCh1y2paSNn4pnq1arcY17Jwk
TcONThg5FFgUHx6kfCyQMAARsy7NkQojPQ06267WLtqxJxPtqbVnCkt9TTJRex/TTQK+U9ubDF0O
ifJ3PZ8WWDDWZ7Tz7OrzwGj2gar6KIcZnbOvX8bxMDmjZHwyul1WiS0fu/FxVn/nDDsMZXGfDbhN
nA/iIv0OMDeoOM2aeyWYs1RCoLlFYPagehVFR48iavVjlU39ZGLmADrtzztsl852eduJ3sLypWKf
WBxz+RYJ8v6HSrMuvsk2wpJ1+9r+Q6tLrkHyadM5sKoaiclD/Xy6JmkZXRhNJiweY81t+i6Es+Pa
VscyMGELrxOOoa8rOGGS7Ncmiax4l2iQ2jOG2fdwvsJZKSvc6QpIrKXkDXL4bX9HhezsE2IH1m6c
0AUQlvHC1R7z81lhry6MO2g1fkmG4DmFWZuP/SrD+ft7Ta9t+UT4c4HhFbocYxwOF2tMs+FG0g7R
rIa0evvKdwuhycZv6flVoMXl92WwgsNo+XeBkjmgRntTfuJIW9NZJi3+mhy/8efEv5aO5Gmg9L73
MhfB1JW95R8sPk34rt9tEOKqSN5qlsow7+WzM3MPliG3/4+QVX392HfJl6W5Ncn+p729CI9cXNuY
m2Exg8jffOGp01L3N2b9eruDAfFyR3RHfs/LRQM/nWrLEV+88PAcyXgGuXIbJ3rtKTPJ2BehSRMr
DLZ8mIXeNaOMlXtJz95JC1HWgwWNkDkdqvgcT8kC+H+7sN8g0qsCPR2vajqb1Wn7d2tMGKX/ZOWu
/y/hRRU3hNu1AsiFMdUYGL3xiiCNoXf55P9yAOEkuEuYe4OcyQo/QfRkhSWiOXWNXEjn31bXGHMJ
lHWvEOazTNRTYXgU7aDBAYID/msjG9tRNGgJTcgL/7N9zTEsLm0WUKEMGIypM6j0ofX+Q8CqvIWu
Q4IrcXKc4wVBmSV8Z6HvTV/zvpcADUCKRbIMAcPSy8erDA9Q2Xgl0p9O/UoLdL0I/fzRUxfT9NgY
2MfkVJuQPoRE8pvW/Iu+BD0j+QAIkXDk3TuqvCSVB3UfRk4m7ATOIE+FuOPIytVd/g3SzD/Mlh0+
+SFpNqsu7uK+VqkBV3Y1B/VCGMS2QCzvIJPUm/OrMuPfcj+2NhQJyPM+gopjA4yyefYhZdQILHTV
igIw4zNgF7BP7q6oM4B0Oihy9sAnOekOmW7B6tLfi0Rmjypp1ID6qIf4EsjoF3AHa2ydJ9Aiu7XT
L9QvHySNSa4ZndG4mO6HB92VaxXJRNY8L8WiyhR8qPtZhF4xLDynCtaRCZNBOb3AFAnoNCc9zjP1
R+WzfjEpEbTtnuYtvPtLKIUul8Kz1bTPLSlQS4CvZaJrNl2IBp14LWqJ+JeqoNrJVXgI+SwBmsuL
tJg9JQWvNw6XYe5Ufdf+gNZkHgg79VW8Ry1TXYcAV7NllhdS0r3zMy3TH98xujz47mcA7S6ZKrnx
Be6HRRx4KhII/rWHUmzNLs5Ps2HFSs7b3oDs4FY0Tz4pahUyyOdHWqzcCDEE67lNb7G7eHmezKG0
P+jlUCVmu7T93QX4ATp/hM5LMgF0yV3nahZLBE4PH5Y+TFALiO2CyaNmuL+wZKo/wGIeRt8VCBgM
qynSP2sk+6WGoHqCp81Su95S1aKJJmUSw6tWOssLOZU14x0tFk+4JfX9zv0fxPmbaczm3D3+JnCj
nYM8Uh04FUCkTbemqttR4z8ENncA2jYB6xnquI4YBdarn73bvkCKZfx7uioMujW0rsqjQLu6YKD+
84Ci6Ywk1cO3SOEirW+DY+/HSiw6298dGAUGQbyNBXplDmHjgfu9R1kmGNgkG8ibqjn3eJF6a8Qx
TOCJ5/g695yfgUQKrlAX0lnCcrZThAhi2Iwv8iZ3fAoFdTKpIxHsv9JPGcVaryQ89jGLwy8F3YzW
hr5UF+NGv0w3kzQRMFcqF8SaK08lTvNtwQqZPVPaFQ7CqDTSb+lKY9YaUN+g16tpntcUhyikIl6S
4a9okkUUM4BmUicxAdPVwV+dFg9TySMlSzB5O+I4e3qiuA2e9zx11xrZoSFTSzD9PYUg2nMKPPch
ePneeZZ9MXVRarGjOHuftrZmmPBk/0z1uR70I3MplbG/QFuwOVcd1a8Tqkf5P2PyMxt+lC8Yn4XL
25OXdEP+xjf5meSM8FoctSb5G5zS4tYGe06UQT1GMnkvOXaSAj1H803n7olBwn0oGfWlj0kP0PNx
dXUcYbR00CoATK8qkUjQlkeT1gonmOHHwzctEyyt0q0+t8jiWX2U1k2rD3U6PkD9uwj3gb/YporJ
rrFEngDlHlvfapOJ9yGmX4GJzcrdPB33NZ7nBNR2EbnlcPRENB/YMPGqh3Xlu7tf0LXiq7xonoUB
WwZVjWPykDJyzGzdE95UEgtr31sMZsyW4Vaqhy3MUQrLzJglAZRE6czipkIUMzibxw31UbwgEA8z
Rh96XG/61YKeUk39gFKpHXrFTIRocDm0sGQYpm1A5zhe99PuNHgWcgSu6dndrjGQiPyuZXBO7GsH
jGMcptPNkojd/VClpgtMsx9n8MGTvJN0iGiIdEELgoMiGMqPLTm8ZsmJM1jSBYLeOu9dGb0tqM14
FCTOEU5nhhM5Yln8oXVNCW25jDzmRG4XZKBTVBoUwdsXanQIvu0wuorJXxlyZY2s6+Fs+W7/cpzK
Dbf2IpsPu/ACIIl4/WMDDRqcCDbdi1mc4CtqdJNeO8SIsUFW5TAL4bU6XT8GTCwfizFUwN6p6YIw
oj/q1pdZsZPknGScqtaVQimcgbMRLfZa1HJ3hCKj8HyXBb9HZhTzBQlYdpzqNMvakb8iYtZaovAi
JlTDG5+YTtugkcZKKU70hRqmAl1KqCgXU6dqHsOJis1HiYSdkhFXB+jeKtUV/qBpD00srdaDsSlF
VAEs4recb3HMkGLp76Ulv42dXIhPdD8v3/Dzkyv6sTro5NPlO23vKI12ujfMMPXy7+YLdydfelcI
L3bVS6sxnP5sMGXbjNvXBviacCvJedHinAHA3vLBZqUEliJd/sq/1khYsNLBsYxa2W4MTxPUi0VJ
bncWFGXQHzlN/VFw4ZTB8uWbSctrXWWRrqMA0PaCTV+tLASW0BBR9N2rZllPkXrkg+sSNa2GuVoW
ki1FiMqklPcpSupcVI5qAFi+wPxSn9RwmoSiCiluq0+cse5TUvO2ccK9vadlVS8gog8Qo1LzPk3M
b6Qe0XLND9/itY8VkTfXcsjWZJBfN3wlqsK+0MDz+4GKb0+ScR6ajUk8b9ilY91TsKVrow1DposR
FQef6OdB0HIWnF+trgbpHoToIq6CWHGqDL+3NHqNKiBfdv5NKvbAkE7xrI+FOe+MpNoIlWPflHGP
iAACU+Gmi2+lgBhn5u9kB+KxTKUYUFK8gJsvM9bk0RL60Vu1mCrmGu++llLZnWaYBSLiEgBbFyWf
Yv3dJi1l4QfvS3koHlQ5xtrf2zm3E3FyWD36DnWCBvGbXfAUmxoRt3f0kIeV6jh2xKrcuzQLhMmZ
CCtDwUAGZvfvS/HFzBRsdvTsSZf7HvMT4OSmRShlB0To+pDrNRzPTJksRcLmi5Mz81GefvGC8AVX
q3wdjOc9cp9B+x00CU7MZxE4G1vZ2f2iSOntlIpNvfHYiNbXItV1udS98c/baKNRzrqw5y5osL32
lIRE+hxu3HQ9WJUmgFn7yICyU6QfcORTt7GUW7Il6tOfUv9uhEvFuKcX/JeA+fOt8xAMJpXJ2GJ1
1YUJxiPJ7H57AO2rtu4ev5B078OeJltLDu/DIwOIp49iK4mHJqrHBSBgKgx1E8fujEqkq1uT+uj2
sS1NGD3FLKQ+0W/PBxhxFmPV91NdtGEMQ35Kh5UhMotz4zNix6A+mHVIz5uxl1VKLa0VaiHbmTWP
jbSqKEl+IO2JjDaJq52FnWTCg3+1/QN8xugeomqDPKj1myuhWrv+zbAxuBxOviBgw60F7S+Qx98Q
MYuAiV4lxI/T/Bk5P/Hq/qrfg7AUHssqJdcuM+7Ft5pTYEQSfMat3/s8XTXX8zaw6Z40AAlEn9UW
bBh5qzlZjKXKFduPvRBQE7La5DLxRyWMORRnOlXzAmd7fmyENAa4atbcPSZRW4EbSW3/61Vg//gE
pUQA6M4rtCAKsMqJ8X1fVuERaEJNh/myQPNgJRRCpbOXMqX2pZaj3W3G5LRBoCOAGWYwoC7ea8XV
H5a6pE2K1wO3DVkHTzgjSV+27TR+sBVmCDqwMxocTyGHmdo/qOmgVB48lFFHTW3PLmJ19UBFGhlz
iX8B4MIUFjtQEYY7yzB9HSSMc6k1qCxu7yly6zj0LYCfHuJ4pa2wpO0p0rMvwbXVgGsmJiDyb2Wj
/M4Bo0Nf81/+4MsUchzak/irMSiEsBXA5h3iAdtVNj9CDOoh6MGDN6D8Qw5LrxfpM7xwLGGUFdAP
8XIakjY7WnOF3YUTXGn+G01JstYY/pFfa/mQCUs9/qzLxl5VYBDVQ6nf8aEE71WzDysDpMOTfg0z
Wcthg0v2BsNxGYIh81hjqRfyyzWmuc+dVwiJYkv0IY2gQYZmn1G1AsItx3r97zWWEXTQLgPcdDnF
DUVtlWmGsNeLR/G0qDD/1pXl7UXxaqh1QdAUSl8oZB/WLyaNa4icWYE4QRJ6Qk5VDYi2y76cRYhQ
ax4Cx/Yr470yjhOUt2sfq4QVeiOHLITcVUilQvBwjfE5dWdaeUcgxsJMUJPUY6gNCAZD3iCKG4pX
+RUjle96/rtDEfbFyDt7j+nwLaDJyy44gz0WWX9ADlBITu2gKsnDPEc9kujFDgLtdz7x5z6C+WmK
vXyB7xQ9SCk7c3WGPbdxnpTfnrltbeEVLho0JzWPSiIwQg8VbVQjLQjKq/VdHSPbiHxNgeMIWoM+
veY0fGmqq8QI4V8iqv0lVtt1Hs8PChD58Xkbv9sbmCNNGfKcsW5b0b8dYeY2QgGw3coDA+hx8Wv/
L88wtyErvZy84ua5wxw86NGOunS1LLRw/DmysNu1ihOUEZ1MaQXCqFsQXYknT9wiMKhmKG0VBCFf
Dy3+Vu4XW0fo+Bl70OMffMfwRoUM+tj1qCv0N4mTFPnPogiGtdae8UASCF9J0UC1Cj9Tpek9Lrkk
bfF5bsdSx6UP5GDK/rMC9s/vOSg4XinINoS8Y+2m4E5T8c8pjVcGm7bfEEW1l/qnb7gVChyFidYI
5+2vEN9uq8iUuMHtaoa8W1CzQI+bTuU/w1TddZQS703AYHGo6Jzl6IUKbUQyzdLkc5miPROTas6u
TGa9+Ma9nCoVnAHUNGZTRt9jJzund6NUoIhdwKngYblgab7y3SWYfK8vrS9mPeJ2Xa/qou4MHH+I
NJqq8/VEdH4Bi0/Hrt869h13Ybp6UBUaby99RQx6/3uvaznLR3PDNMHiL3VLz7efW/ZVFRC076s8
osg1gxZgw9owHLGglg1wpSf0dgR3o1baaEBJZRQ6KK/83DXTuwYiZhYB8jXg/G/gCGv45PCbB9vq
u/+UbOX4fx20p+GRZhdJGKGD72f408aQseML33nfERb/ZGbMSBdmAPRdxZMHUiWSnD+CCl0xNgEv
JTFX7jCkAfDalulN9zHQnFjg5KM/jzJEfB/fQAHH28P58SkuFgs+N51SvtAZaG5xmPg4AX1ztc7E
Y/oCELeqgPP9R23sDpS9xrel/0+qQNVqBLl98a3ORLGdCPEZBzQ46TLu+lhPhHLuYOyocetJILRv
n+763X3tgVzfIzPePUNCZ3CV9/LblcFhxaLAo0zB4DANflYtADOBrOhDQDDS1/9SFhRAViXgBZUg
k0Meg62sQb9GK7An9Tx8zS2k33fti/6JhD5FNtvvQElpF+jFDm54t3+uvHuCM27q4R4hQcmUuE4t
n+A2GARzH5kq5LemQir0NPNahOA2Ow15EcXD0LKH4dgeaGhpX7wynKyGwSXmxhU6ppCod3/zVNqh
IRxt6rogzfOBneORDBbGJ2mdFrXupi8GCyLe5GLETiG3FqC6BqlcMoJZaefCTltZNxrYwC9s/JFQ
Yb628ky9UY3LEGONhy6Apq7B+oKixkgwV9SdaYLKy4idwnDuw+ejDL0mteWVJ2E2WsdS3bBc3IW4
LPzi/NzC8qm3RB0IMeYhRNScQMfqFXQdh4ARHjFzVFd7Gq9nH0yLDKavuRENLF8Z6jhTYjFbNY28
d2JUODQ32DiM/ThMxHODV2A6peIyOLeD4VIZih2IXh80prj8kZrUVyTnxfQiq3F/nd7rfZ0ILd4M
nKfUbVxs4l0KfYJwLdcEDku6qfCmjLRdguQSy5JdjwmCyWTElp7zP+rXJgBzYk1+Aa3kU4K1gWsi
OuNP6bhtimPSXuBJCtcGOWbJ0P1gxyUZQK0LBNUkBspIr9Yeiin+RfQz4nqnxjvrBvzPVIsvVlne
DMP1Ql3xMCDoypjom1jY7xyeCOYG7REHaDjAsxqWExeoueyl9EUpbKG8mgeBfqibcj11rGb9N4tG
aIDcaB6ZGgq2iCbcM0A6YPUiLNQCrR3I0/pD5oQj/+qPePCZdV695FuA93gBjHAebyGc4V27ZMeT
WpFOuWcrLwoCFwsnzWJWQSQOK+2dbCyPt2GSJqxFhMp/9Ksks0elauOmau/F7VmS4zsdiuwT7Nun
qX2NkMUavlVZf4/JjCNJz+EuOGhnZZ6oIggjosl1tCU4GNphaiGZlZBJuM648CSLkq2/KkWYVA7q
lnqxrKuLU4YBRYzeJV0TmW1ZTF/XTso9pN28DQEJZ1rdxDA1hikZG4zNiGWhsTJD946FtgrNBSGn
6jnU9JwZT/hTPFVlva1iymKnmfs84Cfc0OZCEUd7td1uPBp5lsc83wiCCkTj10uBe3s7Nj9mgaCD
kfFWp+7PkEnCdsmSAejTvCqsqkD2xRstLjHV2E7C9ozXeV3JGaeREhoVIzcsEbUacoIej+Czx7ny
YWSuc/4jarSZVG9ubLD/jdioW8iT+1wDb85sdBEktd6bJZhfYj+me/PnOUghY9NauNO0vjjedC37
va6HKZmu5wz+LdRImqSyRtv+AyYVP40a45cUML/G+W03kTOtR5kPXQwZ1gi5SiSEF651A2wpn6X2
JhYz/AmSpA4IaK4A9uwb3Xl7QY7ydgzChxBeXxJ01h5AAJi1YDG90QyfetR2bH7pcOhvlhq5QHe8
QGjqaSzkB908+tLidjb1kpjzMSa4CysNd9AvMND0kDgMSnTDEeqwT9yyCAhD4JogA4R1iy9vEjt8
7hPGJueQcJdZLhQDBRadjib5t/96j/gxNpEQyeN6LKrWQGzaiiZ5Uz8/KZiQcK9QAXIiFVKA+GE3
xOUz07bzGNoR18uGQLr8a2JQKEk73wBbdNL0SWvFRA6FHQLBtcNQasjQCr1qIXVbKaHK1Bz0kERx
oTKOyURL+Dk22kegPBOEQX0jmbpBmy1Ndw+HgyU9respG6qDXwJqR1Cy8G+jfm73T4GyEPu11bmw
wIKWNsxqULv/SxSBSxtTBjsMwwyttrqBKoeVf+/VSXHNghZ4/5SnI3BYruX1jV+m3fSzgFpClIy0
M9xIBL3TwnSiLLn6IxhLHxrLAPQPd9hHYT+aRiFsQXMiMZR7uS5JNQNAdp/+k6+ooebfdHZh1WH3
RSXvg/zqOPg2c+JgieXsom77VsBJkvndlZdz1kF+bVWLYBmzgLHcr+5CAl+EJCvzVN/IeYXTYt4O
o5ij2h69uWD7J/c73VlSX56LnsDR7XecxsDBKQOAjFEomUrZa2P8FyrknqUeeebMyeIzFXz+lrwH
zJeJ4Fb5VPAtbYFJAEOuIgtOsQ+uqaHW+aBGcooOKfeLhzMcpzeTBZQVEcL9phK0EJugPBgNuHUA
bgSYRKDo/QII1pCYvh5jlcRXrBxSrga5oqXLiCpF1oqZ+YY60eF5Y4zaGOePM7yJgemyythOU8Ko
oSCxhE9ptuqC/HDtQfrvL2J6PlGguQcvScU7uL/mjNQOsf7Gcmx5m0r8UktymVMLxmm/Hqfi7SLy
bIZaV2Eyy0tA8i8FWCAh/zzeGnCUZvYZtLuFqN4Gy2Skzr22jngCW5Oo+Bv04XZHdtMw4O3C3Cm7
bO7LxuKfN/8aOw9M8Q7msCqX9uEMYKvG9NeA0TyFr/PJ5ctbayLPmWOpaJjyC6O8CWnbOBQMGtAY
/Nk6I8yMDywc4AHJBtNnVCAUqnEnNVoX627FclsQXI6nDfuhiI0p+V003VO3gSYFARanBotGiYBq
KtHDn9Xf7cDs23trHlhHmzNFn9F6T+1LFKHfQgyQ4bdPOpFqEEgD+yt+pylhrBp+oz/GGe011MK3
R/Bx2khWDyIQAnJb8yMfiaMGUSY4xdmqyL5bHpXOd7BH6nD6o9QDz44jqa0pOArppxbfaWLooF9e
BomotSpNlCfzAO+UcTjVzlGb8PJa8tfAa7gjGSAK3J8eUcQ7kpxDXk8RpGUhq0Q1l6CuQi2ZOP0E
guzDBX9b1UZHbXw/8RZPwU0jM1ZiNKeNWanCOI1LT1IeCG5nhE65q7oPo2zGZaCM+sr2WujU9OJE
szoUPLbWaFK57vlUqmLNqMLl4CKLozkBc4A/A/GW6kH4U86fQCSTAJ/xdasFjOmylIXwlz93m38s
BXjl1LS/dBGs5ep4j+nrYaGBZy9vUKD0k0DfDk6oUJVJJLeJ4riaoH/ensE24iOHx7ayOujToZ+i
82s7zXosKPIY6AViyMBD1daFwZi8VJA0qZGBKndrm8gl5i5mZvyK9shBUlxHY23dPp6tn+OjnqdI
KnJemT0mfgs3/mDqiWXlHpnQaAztsjz0bvhbGVG/nq/WQSMEPNmwUPs40Nhkif26qMa2bx2LThFI
bhuYyLXCuF8gHm+u28ZLizn+VrY4LiNvitMbEQEPp3taZYthLi1WMcsC+bwAVvLPEKq5Y/Ief3gF
KSqRPeO7vJjKZU31UfXm8i8l4UYwYg8fN+M5IPOJF6Sw59V9MkF7Oz7O1B2r4Hi/lThktSnWjJMb
xcbXBngI7bo5Go3QD3vo1W3wDsl5UiEg1YLwgLV40Wq4KCuHwr4jIOKeJvPa4WEGMik0DXJXnI2z
DtKo4iOc3ll59Xy+2IrV2qGXvWGUeGdO/XNFyu8iCyaaq7QxtIh0nayifnX/eqkzDAoEoY17BLiM
D6wdp1O/+PH+ypQHaQuoY3bT+AZKT0ig0xF70AD5cQFlZjpZKifSHKgyspk0TGibbETKf9cR/Upx
ttzIDjvR+265HuRrhWiB4+dxKqjoylXZ03PswrtswJGoUmT+oALe9y4umaRzb0Uny57YAwm1iIfh
faPWM1uXiIZWfn93cKeSFJ+L9Xrn01KhnL6spvktzuUBYTmRXPC9nVFNJsNUQHBN2zpwzgEZ/mif
cZliwIKz3PCyfC9rtog/0IF2Uoz7Kuf0xaHgTw9jZeZlOmtZaZod1lN7Ff2l1ZLvAoPO/2G8/2oI
jWrkiexSa0Vf6q/3pS8J68Dap77NWEFwImbyUf8pUuEzltZf1zTIJZn3ItUDWVyHaCbl0h66o7MC
jBPimgkkIXcv0iZjQphloupew7WIOpu51tjKHAgAx3/mmfaUIL7gh2Eu5oBsDigpcEAPhBzMp07f
Mg1NERxe2g0xIwW3WgV5Gw8N0ZdIMpba6PuAFn9ODQvhnq30WmWVwEW88Vsu4da6V+H2rUEVhjMg
mrED2IOlm8/vwu+QqE816X864ctoJ03+wnI4SK7zTIrJC+1dMrXld3uQzV9dI9GDML/Iq2LloHcJ
A28W2d1LZYvzzM7ocwwXWoSgvGd+KJc0HZnR6lzSS0rBf4wD5geMhY8OFpIED364ceNO4jFkbI0N
RJBmii14Vf8xJZ2Sf663D5sKmNFTL3iq5TnlYvFtOuIFdrNNa7PbKHPVZwkVo0DXzDw+1VfRLXUm
9dfvXuOtvJOdNCsH8IpDYiCBCZTsekhnchu05+ahoeg0uvcXiz9gF1bvkrjpFsogGeOLgySAqZ+x
5pir29KkvA4nDIIgzDesZCzz74NJno5Ash/7lBmMTX9VDOOXLZ0MDIAH4ZyEOk7EhUZy/tFKSid1
7WlzAzgN7iQLdx/bY/fFl1A0evsF8nokmd+NsnkGlIfJdZ0o31FGVpDij9Cr+KHLzC1/3ZngUiiv
Y95vhlxsWc62wJMPqq4j24C1fZ9+iuv68QmROwrwa7tgYcdhf4ImsIIycqEz43jdykzyz3+rRJDB
hmA0/Y8XC5+2Uo5GzG2jrl7k0Mn13XVpOoixeb+z+CopNUilFNc7zHDZf2u7SpixnsfjApCBx74F
a3kLXqa1e64aYfTrxgVpNpTIEIw/04Yjo68O6rqjRmxP3CTRl50N5+BhNjLvSKLXtRqoKnDeD3na
ZIHf1e6doTxTqsXVCOq8Xn4W9hTeV9pX+HiUq3gw8k0/Ya4btZb2bGbbuWbTtgjkT/yWt7Rt6VLG
nx0O7P/VV2Qkr+Z5lmHphrADhN+VkvvxIeSK6kNscQ6Z3W/o+92ZsfwK54F6INR8souNIGunCWVd
lc1g7H858tPClmSJpfUqF1Lb2KiCivEiyM1K+dMNbQHysHcd+pF1o2cfC+beRp5EEESLMDSOgmuO
mz2yA81sF4n6FOWu+7TgCbyIP4/EMTq7DuAFilJy2vSqlQku8JgwC+E4PHeLXYbYUY/dqJ5cUZIr
ACzU9wf4/NDS+uzwT2rnMWCM+CEdgOyoKVtHvUuwqoRh0hICageM9C12zXb4JKW4k+GKoXLav4U1
2mKBHbUPbIZE2LNFZr79JwQTl5k9Jp9v+Dwi/H1dNxR//jYke6XlyXjIX6q7X3+Ga+obl0ukflg0
Uz4thMdj3lUgt90xp9SWWz/9blwtaToVd97XZLRL8tIKITDg6YA9yA0bJavq4FS/SCmSGmb/aYWT
kvWjVb1xRls5jbBzuwcOgszUK5VwSGWO8+By7VVRcRGAGbfSqwJoNeJQz21aqxaG5m0R+Vda7qnM
vg/Sx1x+jyIyuS7SYmWLg6MQbJtLQUraYCGPu4UYvMvfsIAsWAymNG9xO4CPjMjWaY+55RywtRct
X6H2lqmKHZWKgeIHpdfkYJMH3Dygx0qxlA2bz5yQDboLQBio9Nora9XndfP1Shc5OfaQvP0VEeAa
DmDC5bLCFvmPoxnEAkwP41nXSSXGyor48gEYuDjsFoJAyZEujXTN87IzmXW4lRMqWIgZ12VwTwsU
MffjWx1YSQWu+EF83T4HwYzR4hHRDVaIw5bOxhdmGpnC/cukJfa/IiLVvIYvwREAG19g13eDQa83
ZXB//2KkpTK336wPmhTAhOGAtA1wINMYd1RTTBdkd9otqFVRbn85iZcUDlXvU2qweJ8ygwwpVWeo
xOSkGyVclmAxagG8f0ZcbGFrjPpvDZ9Bo017Ko3CGAK36whKLdxTaXJSZrcWovV2B5jUjrMIM7fZ
kB1vOOI6R35GjdLnhybzfE+oXKgdBfPvBSE/mtMS04L8xU2ZrsbYCEcHeeCKa8wLQHlZbb5d/QgC
zydwT7HfGe0Rn+kDcbjE50aXD4QdGCrnmS7Wv5zoYOzcnDMVy32SaMsNNZHNvvETNRB8Zn75fDmE
abLgpD5QQbwrBljiH8wXapf0XrEHrSCLFgNt4WAApXy6fgb8OmWKoBePYzBDMkhs/JSyPsUwWaHk
YFVhn4fGIzXYgj5/pyr/KD0R3ODHPwyXZlJDgXhbk6qpc3Glr2vrtH9Zo9i7eESG99StFrFDiPT4
CvdkDwFGtXNNFBI+qZHq7m3ciXzeiusv2EJQDIztWvvjcPWc7daoMan8aUrDwPozQ0Pvo/tBgMHi
Z5vrX9uW1CZHz9rCxTs1hWpp4/It3I7iWHMR7jmQq7GWDAJXTqDsvnJf9bRzI4KcfhfXaPmXagRW
Vg0puw47TDqx/A0+cF46P4AlWfuvl1sNzBirqWUhqIYv5ebpLCWul1LN/85KINLyJhg2Ke6aOo2/
TUi/AzRvMwtZhGb+mDqkX0yHAYmF1oLoVc6BMykFwG1lIqljI6icLoVxxKLYzschdj6PNqFRelcd
Uobgj0dz+FA7Mi7uinhfLsrGVGJI1qcO/SR2tVFjMf0aXBLvwhOndXgs0q+4+dXGrm+ZBU/fMqr2
MXnl8ZgdRubUKTqLlGixqNyPBuE1OXzDc3GtghNrcCT4/AwMJKc1MDRZOvpqmogq4tOTwF1Qqa3y
yoAzbd42/VieTasPoJScTjQ1wv0HYxS4XRaTu0mg9P2OLYxOpBFIqVSQwnklymShX1TbU4Hm3paP
4ihyIbqK9zKx42JNBqqoEkv39KeFn2w+Vwf2bMkkrAnEyzDo7xdiZGZL949HntM86hSV2IBNi8k0
uUDL/0EJszBCKUTXpmqTJm46AmsynJEJY8C6/fINgG0rgAKZ9vmQPRLrNVs0fsZC63ZJOs6iiht5
xWgu5ok4YpNRRDhkmuybfkzBrUizDY07xgTTN3iiHKdOOIxip07BUklkr03GP/wdLYyxDlnDA6h8
0YHWaeRHYGa3e0OyLJVDcE/p4FCoTOfK37HmwhO+OsyFWO4wOrpJrXwyJAtHStYot9lxucnuPtts
re+/y/SAuR/dvrFOV6zTEV2aZF+X3XhFwazKnYP7JMDZB/jZrHsjsgGSatc0H4PHfS+Av3PukU57
lZbNocDTGZ26ylNwI3Ow786uip6UFnrsaqzoi0hmEeg2tflrZZdKLxYv6bLYtIA7bEdvoMqY7Cp1
B4oC0QIvYPK0OKGXJ+kSbmM8dmWhS7pWZgFfs4ed7yD2s2hCCSfXkWWSNA/PlHGv6NpgCJH+GzAM
TIWljQAJc0Jc1v3cxvEmVHEgWkN9Y/Hqk+OOAwf3q3yXpSBB1uAKdzL0vCcDbYLOwIzBj5dwIdMx
aI4MV2nhDND9nmIzmpX3bxCM9k5f3ZyEdgdvMdi+zdnD/rRC7XaxhaTyBSWhCT4Djko7PexQW6p9
xpRKEVEdPi98t7YBOFWtw+IZS0HgBHqnordfDqbzDnrnUQMW8nWiz0J146iD1f1w3ecAMhjI8xg1
MaVcD02QnR+n2SDf3E/kdsBJ0TkSbIkKzCdXFGqIpS4X4xoX7WJ6WRFfrGPAiTnaD+xBKFxxeSTb
xFJLi843JFVUCmWdMeVUYQF/j0wVGLdmn3MivjA13vWkODZ60AOPNP3jQcJDFAwuPsC0aSwsnDG+
VfjqYDf5e2KgH9TkLFzeD4mZFBV9AfBsy5S3PDv2PDobfm4FvqPPwDWV5gf473vqOZ3TjUU/4bYN
uPFudxBbcpPFZ4LTJAeKdAhKPoLn0kFXy13Pj+S8gLQyUSEDJR9K8GRBwTeXMFyspjQNB7c9reYd
6Onb9wHUL0qXoj6RRcOm6LuHNNHRZfT9zWT6ms+DNx/37qHNstGvOnkmMetS/Q25kAx537QGdHAk
Z19R2TYDUxlYO6xqUz+FGL8jF6As8lLh1MJIA4dr//vjwrdpS1g1Ton6wCHH9uvTAobckebDffqb
G5w39EMcLmU+y+AgPiSYYa/6s/tt+9mqwMRCR9GfNAPpXfD2v1YI9rctgL6niBZRegCkwGyNhFRR
Xe6lCeUDoFNPlqG4YJv7ffvvzir4UH6dfBsByYmosTW//6XPKhKD2NOFftU4x7OVzK9Q49QV+nF4
pmakZdxM5jDmKi+A0NAXj3e+gskI/4fUCMuoJFejAx/ZDVnouWWscrPkCK9k/aBctTJghKcCBHes
o0tZ875XE3u3RqwND6q6CmouizNvHYleVRQr3EHMUvOTlfP5j4Mzjnjj+gdE8sxanwCuJ3NQ/n4a
ZljvtPcwIJ31uzDyWC+Jg774e7bBHG6mOpTWLf9ffq4K14T5Uv/6pLbl6jBms3ptY07HzLVcF+4a
RHYX78plH9ybr0l+UVYB9y5JD53YwwFCdAXprs6PTMkIRR15tsQ48Goz4fWBucoxpEUgOES+1Ok/
3WuzNzGg7DgnIffLH1URV419W2WSIXPHSZRIQfdHIhOojGbx6j5oHCAEq9tsnxJQ02W0I3ljrdYD
8KMH59TzusRRBxHH7NZUOIey1GNRY3OY9wU+dIVPCabajxoyuuDtydeeetgg3Emc2f8+dOcU8aBP
EsobsgGO/o43g4dvv+86sP7j4mNG0eMeSIzx/6SE2X4hv0gzKI9O5vdZX6F3rEJDhB9knCgaSNZ2
/ZdGTjIoykqq4395nEmL2AWs/4noa4GD02jWOvRx3+RKBeI3GaZvrnBUfYC9LTQGZHCxNpg6BdjY
akUmsF0Cau/kulVKy0e6w3xTMlIfg9eDXFGa1Ia0eYWhivhlHCseuwXqVJrYoCqcrGscNnieU7HL
DJfl5BuP2JokPtPUBeyOA6sI9izxhJJhru5oxWIue18MWIrBt7dlLI/5tm8RuRW0qA2JSV0epG59
atOnr90M76DaOPleGhOYLumroZ1ctjLHGkiK0eKRqnBpSOhzAVRm7ZmlKA2tFzdJovjLU0RTaqlE
ymSLmVHODdaIS10jGSbsj4fpnG+a4b8srzbNoP7pw4uF/+lOx7vRXiRokWCxwajV97wDiIaTjvuk
ylLZ0zeopiCxvSuVbMkDHHP+JkmJOj0Gwx40wsUagfQhJ0nY1y7UnEfdPvQaOo5W72w9xen/FJlg
gwTjHzQ6AvIasIyMY0NtyIaLm8B/a3iGJuEw8/+TU3HFgvLWhTgpQoKS/lfs7QL9wilzauhcopa/
XTNCoolMyx2gNNeOKNvSH73GQJe2eZjndEpopNtT6DA1ISMHrPr7nm1KovXfrG+5b2JYv/AG3oMh
Vk4o5PP+F7EdYnnVMDt6HOlobLkT9I0LSsHeP45becZUtRXCHKsLHmWqLUS1/0r3rrfxtymkihhp
+i2rs6ViKzW6yYOLBc75S5OJy0o1C0LjQ/SRSh5dyJGcIkFJcJj5Rc+9vPN3FXqx4lr3PQUnZ0mP
iECuvsu4D1L9GTvT1MCUJmfTyunvut605LBQkd6i82ieSPPl+Z4lsDgRir1G6ToDb491i6ZBFuc0
xxWEFNGj3uAkQTDq/JCYOX069BdADQD4iSGXdWcB3RHb9nNxHIX9+jaAPXNT3Yg+obL/u4KTte/R
U3mDmlW5Ny2VRydOZ2BH2V+yBZU9UbAVGUC7iq9JTFhfTxbS8JctgytfcWbIw4FBzaMczq5h0942
GJvH5+g0LZP4LT7AdEr9USlHBnRytYMZC3p6vejSa1l56oHeQUZ4CYtVWo/sLgFMU+IxtoFjPntn
R0WoSrz3DvZkP4qSrIep4mNIxGIRi/T6ZrWcGVOBau5DGlx7Wd5EB7DLL+U3vWHNrrCScsmLzR3t
cFhRD9E4ChKL5DOCgbrERFRVnCtvCDNtAldonD4LdPgCoH4HDU/Yr7yXP8MttJas5JnTd3aB/N4v
WM1z/5oQTdxWyZeuLvLRN6NLDjTc6CiGg0hbMQ+BJLTvuZxx7SoPxfd8s5LSBQJfm32+lzafhJIC
vtGncqqvyboh2nrbHkWkYY81FWmxiIHpoSouFP3Jml4I1nK29Gzh6WqxNAruKheYGFsMrladR8t6
mvSF4H2Z5KxVdVt9RppsElcb3Cb5GZ7kM4Fp2dd/mY7xo6G8mZNal1HvGDDFC75UyOzmnMtd3LK9
b7fPg3Y1SsnMtIyGmX8JSHZxfMBt0pmTyU69N9WvejjbL2E1cBy4CMGnCnYXT61wPFpDWAjIkwFd
I9r0uOOJyVJ63l8mOWOokle5T6LWXerIYJ/BZneaywUkeR78JLwuiZ/aPJEqBbD6tZhNmVQFLPy/
S9hBHRCpTiFNmW5GiezULE7gic+Ds1x1FQVRcR+TsM0bmV3WuaIfhw0K/ot7eozx+iZa12C43BMK
EiOqz7LBR278WYkAoIBPjszs461WdHTvquxcjBKsBwvS08aLZ2q9tVBd1KwToASd83K9O4bQVbRN
hoJUAEsUG31hIVN0ovR9+TN91bhe6q3OTNEAM2joFUnsjcQCchof2gzSXEiunVIu+4Zj8HvhR0Q0
FRPepDopywpCQHud0ktRbRmtkZ+HcoaeQW761tXdeRTQxGVdJy58HM4GZiMLCFE87I2VDglSyPtF
URv2AEoAX2Q2mANvsbV2UHoGdi846+XBuWS81IvDgF5nyF/UA20GGKsT334LN9tdIlMwHE79K8rV
MMmAb5T+Zu4BZIqJXMbQhCAIbGOGpG236acWuORgYCARP3tbaEsjT/Lb8A3/sf6V+MRlUI4o0j+n
o/RxE99/LvdS0lbhnY8h6xMTgU3sWzbQ8BFVp19HAROt9kFhg826h7nAoB6cDImXJjEHWqcOaMXc
5w639Ai5YNcOtkKwcf+BDr96aBybcuqYlpCY4sENYdGHKdLwc+Pgg2Yn8XAEUGSyT1lpx85xcoxX
SnqfCjPFO8kxkH+kAaB9iE6lxTYAbnTnIszWkenjM393rknj5MBVzK8sCOrss5wLLgCwKwzqk+C3
atGtgQkkBlTNO7HnTTyi3a1pdVKqScO8O8Ud2WaPc83Oojt6eQkDlC+uOB2cM0Jp0/kDUGaSiujJ
xplB/HZmno4MTxN5KkLoxxSqcZH1rO+8EjpxzyNYj1ZRVFvbSQ61Dj+aCBN4Q1zKUOtd02lz3ioa
3x2NcuaNKHq0lsnToX1ZZpFCv+FD8sDTYHYUKzGs4/ZjD11WQ1XbXXSaEEH5E39oxpuQ6Ln56QgU
nHUvkTGUxH9frjzVBWHyxaLiAlXD8x4wcoDd5A/NSCv0kOmJW+ShmtNrTSglWQeakHvo8uMJm2e8
cMCs9wksvrsE5IFCEWMrs4s88mC7DBGge7iqpJg783BH4rzN9xzOGXANIs0wY/5oe5aGhXj1v4z1
nripl9fB963KJs6Z6RR7OfhTynfBv5+tGrb7iotj0vd9FBKyWRAJqFloLu6esqSmcfOdfQzt6jgk
uNgITCFGks822DEzrKl+Tz64bdLiEmzm6Eb06Hs+Cp0ryTs77lKmY3GpY6pYTO6Jz97aqbjJoI5Y
N8+4D6AMSjuJLtmDSu3bHQYrQfLRZBXIq/H46nldGj92wm0L2TO27rhIUBiMrUBSLbAsmP0IM8nB
r95yKNRLQ2edUJtyE8bfAfZtRPZ5fqs4/bJh9O/WIW92i7CRBhxVt3OGQt+XjkmEinTe9XFmjf6n
2XzTAmIxp4xm3WmhLwhezXBvRkiuu+YUMmuKDNR6CuAJ6v8n7mEZ6VkkqBvdqrZaYtjJsvuLTX35
fQqnZHWYObUvODkUveQJq+hkgja3AbIgSYGN9sX/8KY3ZxTSFEh9REC8PGJj/jHctI0VjcgYB58x
8+dHzYuBKniy0lQ6OqB8tANxzV9KlIb9/p0ovEMTojNNzDYW3+Vyyyto1s0j6jhUG53yGPVXJC3e
ZBYP7BZgp7dMB0aCpsAp5PAdbuwpJcYA13sWhjsLBEjfdajhT9ScSa4MG3nihSb7GBjxVjjpRQjZ
AoI8A+7x5TD1PdrQ/0+BOBuXcAf/JEWuDWgvr3NKarIVsHinAMzURXX7Jv+sMIgmjKFdABttvs7u
cKxqZbEQInKioXREb9Ti26ytF9QRsBlcrbLT1avcXAdg3LFlazsxDnBC5X9E1kyjeuK0MFaOWcYn
v2JFCRNHoi5fnXOZ7DNML4fUJcW4Ix4Usc1DH8b+M3nEMZHJSMDOl1u6FM9o+MQ/70l+ZmSgjq69
kdzblqfGX8ZT+rk26zytpibcjqxGboEtaaBOgGtJrl6rp+dWqaTFpLm7yyW1P2JD0A8VXzL0VujR
DTFQ8NRMAIUv9OyDIYh42VD25US2QYgZTdG1LkQuOAU/BrTa3knwusfsPcj0BRkGPaCnUmWUZyfL
n/bviB/rzb86ytj3ivpHj4U8P9G3iPQwn5M834fE9qgUtVC2D3KhBLUNS8zf7UtURjN56zp2phIK
Ba3HiPnCLLJfQOUPTB7cyEUpevfkHIhNH0T3eITQ7Z0MnVW/Gvnzze2ytKFnbtIEq+Z1lUz385iJ
h+lojbJlqaPh77gfvK8LLBA7LQsMmlcrx6vRBvtG6zWbsvecJndczOXC00DAJTq/0M+bSDqZUAey
6MYtOErgH1hwbCN2/0vTchL8ZMlJYDp4Smh1h5OcfbDsw/wocBnwrSx42tu2ikdPeSnlOQ0v8DSQ
y4s5DvEgeiCo1gFTMVGCeABFwGWfPxrQoMLTp0gTsKRf9ikt7GnFk+iNTQbNaTx+BKErNaqO7uJF
89DY1ZLdC4qC2hCT+gqFeDWaWw8PkEVCqUf9meMt+CuZ7/eoHo0wCdFIbrm8vsAhJcwUJPlupRAw
TQN3Xoj20SPWC5FbdsXke9hgpT1wzJGcHI9kL4WcjFm4bHz7SoU3blpdSd8LSaTR7+zvHAKHswee
aoj8WPK3eqGc1ixyCA8M6FLnIA6bSTeBnMsAfOtsy8GYP2GCKkbJLn9ManZxI/wuvzuDX0uKkEOw
nedf9MhXitKcBjWpFFlft58P2JQXWjd4NY3hqKXdzMSGe6KWFup7BuiDhoUlr1+VBzznkSocgD9H
pVwOIJx40stP+NS4mYP4Knrj7jK4gIDquPnHJQ4OCDkTFVHCjaHdkf7aDhzXwdAheS2kg0gMkWgz
QxygCLg8RYnWXjq6yUw0QEK4vOnkoFDqC37B9oNrj2tTXXhlfkfllCiZdkrEmH+qJ0CM5UC5rtvJ
kBmuGh+Scdv8I8mvJff+2RfzTLSZS7hAoTvagjmougJwSzgClGfATn1j3v0cfEIKPT3VemcR/KnA
spDsJAjc/MtKSybWj31chb8rhaSVgziSWFcZbM+eI/XUc/1mq0BNIX1v6afy/TcNIa4lMQCD6N06
Y03ZDtQ71dsEZWxsVXVfMcqzDCJfvjMrQLTOts/Y9E7IXtGYYGh81hg+h5EvZhmJZ/esH5hpPsZs
ayJyN/jFNv2fiXsG2tJoQv5YJ5WF1YUXnfW5CsdoQfFZGBjGl/hcN95gI6B7bownv6UdIlqiy8ja
wgJl9zdhWD0ZDveHsLNhvIygd5WZj420inJ1swqGNERuFkfLhW1KIyk39QdSC/uzoS+RGXWl1lhU
Cqgb+WBMj4oRxc1/YqHnOlHWhFnKgnQHzYU31Sc65AM9FJv0PkPhMRnqLLjWtUCOK3bfL8jiDRZ+
kKjayGkMPKUKa9pPy39VoptkQWafcM/Y2NPfnxnyFFe6dreFp445Itx+UmqDmpYp0S0l7vAPJgpm
oI2JZLPILWKzmBQhyahzd/rC5jQcWtbWRxz4xLuRlIhhZugkJcl4WmXw/n5XiAOap0fXaf/4kRQd
Mzd8U2utWR0aDRdBDZTLnbCE/50xvPvDRNBnxT4R2mmzUNNzGBhHl4k+vAg1Yr3+IDgaK3ZtWxB/
4pRWGAp1ZMed7HS6UHm04JHhJPD2ef0Z4BQ0djJPiXsJJg8r+f/2skSIUPYcGx8iQhZ+dtMpRgwP
VFh81QNYhbCE4hflBvLBcDS0pWKomG8cwXQqYxZwi+7GnCwRRfqq2xxaGAE6iW36Mukfr0S7KRpt
71JrzBb553Cbpu6rvXixqubZ9BNuRFLL+dvKyP6gj862mAyAftIZiUvaJzGOFPGDIGFsLJNkNvuV
TKH+CPH/DTY3l8354g7C1EaitxIt95FE94AuGlJLgLdFV59jk+ZGkEXFCP97cS8SCLnBEFKOy6pC
6b2yzyASg7HyS5f2URA3ryBYVoX08uWLt7D7BpWrg7r7Zyi64WTeMH6zT2ktn4FDkOd/ciJKhMEA
Dmg4zVqTzdZbHEkImdhNgdeQ/Uy4ZvAk4jVvcGR9O9x4T6QuHmQb9s19ofGuf0rmbVg/eVc4VfJv
tbH2Qc6Atcv8ovtIGLUcPoIKw/T8wS8r3nfQ92hrnnFa/kagMyIawuyO2YDQWeT6MaJTY055mS2i
JF4XhSVwpmtRswll0ie0FAfpEMut5mrDZtOlZMDYSwKRA1zMbOKZTH8fFmZ6pwNAJijdAApS1asm
Gpicsv73KC98shQpBjyGaoUDF1PSSjYKkz8u21pP41tucF11ivuXok/zg8xgVy4nqvsrs4am0m6h
LV8DS9BZVnYvlCphYK3Tbs2qT6Ha64CSoz73CFVN3r15j4ClKWhrSmB/U7A4DY21unUjAsDflk7D
1Ku2FcAcd/+XJ1Rpb54XxvTRY34d1uCDHPcPAVS7NwsXbgU8gXUn4XW8pTNgAUGcabnGqZz9c/yy
NzAoYVXQshJd0EADpQkwiVs7RUU9GLo+3tVdRtVxPURnJw3LgV+F9zmrFTsaodE1IR7d+ByTMtFx
c4vyqVgtUu5Elq050mvm7NicBJai+QXo6jvKGI4xZ1vvwRisxHsS+b771YgJLVEnVfCxjf6n2Dul
vHWhwTsy0LREuog2KNQ1NaJlbesg6lNpyFasT2va+QUt8q0tYeTc3wUYBD7KOw4VWdf9/G1c0Mqq
OA5D7P+zCG1MlPICZ2Tjo7E9fG0L83BMkctCR+p0oMcCR8QaSG6i/Rw3zcir4JiKr06NrCt7spH6
tIXnjkT7Wuwg9wK9b+ov08Fiapo86GxKMJsiXfbdUvMhlX+o1W3l3ipgG3AjyJDC8dFNGGI+5tK5
VhWSZ4tpr5r9gccmsdDetH3VUP78LdnuO45dwgGRRXbr2W2NctqFvnICbClp+dd5SLGsMEPc/8ji
bp/QX1lFqWyAtNt+caDMwMhWmHhqhkDTlyRMOiLgg1p1EcHG+UX54dZbmDZ3rDdXGJRb2qR52Jjd
/A+LnBiUKkeMDWOhLZsap8qFbVyH19L/6P5tjjQ2yuSNapea3LKygWfMgojPDwi9GSu+Zs4kwoPq
vaqLHFX4QDMj4Egn1XqUlLOzeYPZhoEEFTr9F3NvyPUEB9zYVmbc+6aTgI3ek5Lbbo8JRGHfCD90
GAPmlTTO/5WdGoRkGjwYoKO9fkB79UhzBCbCjNk0BvdOeOXNO+FopIp6e79ShmHss7boALqeaRjK
CvpBPevgOgZNo5mRU9uAH+mVNjhySiDhRlkREScsBPFsvV9xBycrne0gzUWNM6KYiwdDTPb5fsk6
lhxOTaYFnG8Hkpb1oPYWvhSc8YIZzyQw+CMRcNvmVUuJcUWVEPTvYqUBZ+trbEFEM7UVrl9IB2lG
Xc4yZKfbjobsPrG0a9faUYldcSla0RVVJdoUVBbHpZRe8tJXbmVo8flYQLqRMMOR3cudVoZ2BAr9
PJ1lv/vM/G+KLVPM3lp1TA5D0mSPtnzLMazQWD7DpsHEOsn9r62VVGgyJ/0VU3RKkvvPOXQNj7/x
immfJvIU6FY2wSljYCY4n15h7w8JWY7MyJN9V4S64pJ+az2LJ3T34Er529ehsIZzj+BavvaYZ6Xb
AG/84bpzY+fBAKJi+Aa7Ip6m4LTS/AZPLKjKr1hBy62cuINoy76yyLW2mQQr7hllakn4IKKcN5Y4
/VFsPmwiqQVc79CYVB6QkrWPicunFthimk7J+yAVOkzPp54eUZ876T0glbe5xajTxzDjMR7+fHYk
7rGJe4DDtM1+4v1PO68Tb7cXz0xJXeWfOF9XyemfilUcXj4n29u06mllIn+S1pRxMUlbV6bbGhVJ
8mCSsxNksnd0mFSKcvvdpPIqWnNvBFF4DGPpXEthpHQUlS/933CHEpaYuFTRDYwJN5WAYaQ/R24m
zVtIdfm0Q3Gez6CxASU30a/zjEaO2w7ZeVyeHNAwwlQ73Sb0BeUbQghNzH+dTV6qAkQC0cj9UCxD
RBDXX2/QRL0sS0LnJ/FA4uoXyGFzaAXCF3c7xV4iOW9LcnwdkD5PSmnB+WypIT76+RVDGUiIwLZE
XzJl7pzMrWELCdbT83FpRBfkf8q5CZxUcM9VgX/Xet8PlvpEfHS8FC7hSEnk6Y33rrouIDIe4cej
Rn7rXyhT6+62rLYa0SP05nhS7aXCkqgEzzwRk8si9oCnYE4sHU5BrqWIw/7od6Un3Ve6MWgN58IV
qI6nCVNH8aHa7smmGqMPcKh4wpOAaBjpTxlulGH0lCzSF2Fwx9oacmAJV8gK0LENE7DTJTEYpX1g
U5VWz+j+RlNXbIoyGEW19cdL3FxmPniMHj18Xtnw5DFgaY1K6PaPoZkL8M5Eg61OhTfE68sp60vS
ms7cKkkHHXz101lARR7mFm2vzyM4mARYgSXFXkIXIgtrcH2mSP1gAZkETvd1ggrlHLGqFnDNMSAC
0OxmIykSN3hXBw7xvC+XOMheVlmY+5c6t6rSYG+pd9RfD0gMk+EAeSUKfarVASkcPXvPHGl7CBcq
+33Ew2JidzT/nyk3VChQSx0kVdQM7jJhBpAbT5W93ZKd/IkIRbZAZOKV0DTeFOLVO+ilcKCcnpKj
6104iOEWGA1ifkv6+7+lyRyrpJH0OQXuO7FOvJv+5yW845egnxChbTSJUYJxUHQjPmXijQD5edTQ
kfJq3Aqd9giBCbop61NKtyqshC1S2IRgin2lc0HJQCnkVgtzjce19gNo1o1uMMSShT6TIhwt/pTS
gI8H1M4fmAHHYMNxejLX8Pz0I2G4vi5MyU+5pK2pdwLLNZ2z2M9cDqh2MXprJoxVt5UovLDPIDfb
N02qByHEDFjcLfXsrHd90GNrn831L9wf+Qb5g3+R/qZJ2xWENMAd3Is8/lWxxN6114MiwHii4mTR
QBz/8pS0WfVUjc/R3BKF/C2w7N7FnIW4cH8+MDOBvtsKc28gC7F7ioLrIbqAtgj8u3Y/7dOKsP/g
QlXDQg6ANMmVdyBufyW+VutuZJRkmw2hwHfOcaV8IK8SKxGxF4yIy92T7sD/0vNumIStyhMlInRC
tF1Bd2zAG8W+r0B4A6UKoJXNvSB4/gA0KZHLOwwBawIS86xMMX9wYiLwj9m6VAAYj/ZkZoBS7NV7
MMCSIgM1k1evRRTKQtgZ8TY5HPEN6vgnAKx+JydZWQWZyn8Iyhg/lmxv+t/WmH75zELjFfL/pY61
majOyLbAbVshED1wryYFRc3jCr/wTpPtenmtaPV43y0BgvdebBp4iJMACjqgWGwuqp+LHPCK6LIA
jBwB2q9MUUJ+QRsHda3wY2V50c/hKR/tF7Z+UJfSNIubrx5U8YF3LsJxzt0FcwGdkTagGxus0qFi
H7zDE4x4YBGMvyIxstu2Tt/m2grSJ/ufa0QNJXnTMSrDCxd6r7/4htEvzwfD3Lu/mn3ZvDkxVTME
dgzZwAaBUHTfUbybAcXqApe+pVfPKzuFqUpY03sLAx8dfUYqly7N+ZHaY6oPA9bS6YXqx1VHzb2x
1g9gFsBkHbX3Kf6jgAdNSWRGVgwqfWQ97Zcyqu3LmF/HmVXKt65k5Hr2LW5flx3zeYct64ieI3vf
ZtxTL8P7zUrfikZC+o2H9oN5IW68j6SxBZSJJrLtWfJYlWRvBXB84ZSUTLfNN4lEa3ZjW2n3Ct0O
oZjtBkW65RuEsw7WdTWC8aeEG5nAB1Fua4vB6sZl0gSsP4zvQPOHPS1CFBLvxdjUNx6SvFhTa+QL
QQmHn/l3g/i1NgsY2rgWZsKHG4QV4+YhDG99CLEbXiftF/iN+BCdroNgrfQp7hoTLqPZtgX1uv9E
0I1Pfy0wzedzI0VzAmXSuDK0BFliDjAryh/8GS2z06m6G9jFjK2W5FmLSOUqIGe84I2yNJq2cor8
mNlKtBSRyUTxtYnERZ5SHEhSGTu3AD29IBwp3RJGTei2b+eeA7sv3ZnRYgQCmech6CddYtnhgtqZ
BYHSTAHL980dZDpI2txC4zhegf8Mfhin1ksyowNetmpjnO3mKE4ZQZClK6LUWPAJkopDbyoAyttE
IwTQbas7+7nnk0Pi4R0YjICRXsUZUiVw4aidOIRT9dGpGDz+BJB4MzBJsz2nbhB76CASiOh5dmZx
5QKuC9kKFS7B3Hg7A2LIUvZ1D7LtF8nYxuBj2we0/y31dP5ThNlskU5w2TOK5pGv4aO+bUlbWN37
B65eQTxzR2Om58qqo0sZ9joJi4/MibfLK6ZFzoFACNbdCuF9klY9VMfwMZnR09voOQ6/YJzYaIhn
EmceYlH4TCMI0kjHX6+WFJbpH9PI0mI1rSMAM7qXBMRBPjQ1SJ+GPs8Zk3IOd+dY+op6T1g7Zb69
Lt09LUlpHS+ZnxpL4ExvvVt/hv9ErX/nsK7vK7qD87FI5P/9NKwDT68v2XzE1Ln0l2ALhkrP/Rl6
EbeiAMKh5FLCH0ytW3DCEYkc0zdpcPte2r9qCCUzCW3q4fvUkorimCxBr1H1BsUVzftImLl80Gdf
9y5V7GctD9Eb7VT2z3JUznUv92j8s/13y2loJWX218ym2w4AQQ42m1+tFH9IMvW2fEdQLgFTbMxm
fCQ5l7FA9seopbWpFK0oZ7Sd2k4wG+xgT/ZnHtOL6Q1sEsnaiwdOZgwbHn1k6XqgfFm8AcZjJMug
6swxg/hCQPyjhqksxWKl0iXn6mgifXg4HtfXNXlbjEcyJ+2ovBBFx+FrOFiN0+uN18rg8eVc/uVF
zVssX5QuyBu3QTKET2N5ze/FGqdtgIQ2BFJep+Jdz9H2PyX4xgj716IVeviCUG3+Ub+ovMkmVYiw
7pLy++bUUrqZXwk4hIWi45YEmAMVYn04jhrYvuGzDdx5uCQ1t6wfOGNYZdy1yDbNMJmIYun7LLER
JPdDRuLcLduhKnyWnJSpA5hliRpAaLZy1ZZVmykkUNBJ4v6m9WW663/YwUO0s4XgswR53trRI4jP
OPXGBIWOWuFP4wvXgK70xlAwvilFmZZeYLSBvijg1eCiAoQla413aTrpjs1ChTB32MsgiO8UZQd/
PVIFWg8T5Rg5PDTMK4jRrvfXv+HaGflT6uQlETymdVinsY37k4x5R/utCi2BU3gaIVth3ZPW94kY
GypRdSB74VJocKCq0xk221SJ0LCAMhFxlf3Su7klpTT1YOoHcYN6V28pwpADtac1wtt4faWOx1nq
vMot6scro+2/d8aWGF5nrhVwnSjr7+XJCS997CzgMNUwzWUM6YQ8hdZPUN+ZU10Mqjb50ES71/qi
3RD3ysFjVl2kB4hzN5uPBGSQFnZ2TttBPG8iAXiHaybmupTMSSm5FG0zaIQwSHVSOoa6Q+8C2tVg
5/1YvtlQnoIC5WJUavDnLzYykKbKFzJQHE/Rw6qzZ3ebg4B8BmPMHWS8AHQo4jMkl5SOT1xAVTNp
ZtJn8sMC5PWgnyOpgtm9NDHq4aGgfkSdY47fetIuBTb+SedTptQ6FEk3lHl9lfERwOnvoTg3h/wv
n7PL/PR/TkXz4mR3GdSkgXN/jeQxDNA79Mtmr0agzElo5ni/xYF7nXxt1iTMYC6CA/5se6RAUvmA
3swU0pR20ATZ76RfbpzplYWw27JpoBtP/vrt165x5SeT/tE/UMHOSvLNmfSyFghELXUnMUNrZGEn
aQiJGCwDmx6xKI0TZGWx5BVgd+qzTxKZnroej63HmOwe351l+2NUFRQxG+tGxtJBVrT02Awiawp/
+w7gD2skjUZeVelqNsa1QDuJY1wh6NKmeD8aucYN+G0EcFj4AVcrFRRTA0G2QcQB/uf52jMsWrTV
crlXcCJK8Wt/qeGAu4B+UQMxy9iuPitDs0rhpDV8X8dbnD989xv+lxYJ6bDpeU0/Es/r1ViAAZAL
vPvSfhg3CJlZ7M7nzKuBe6K/Ie8jV58SpNNKwd2zTulSYee78nlzEzXfvKqM9bRM60W+Zd1a1YI5
xLZPEhX7V1YlqHOt8KFKJpOzeoLxrET1kolPilzkD4OGOw2buRacDF1NZ3cpJ5FjscLUwslEkB7+
fZD79ccKyVLeeW3Al5ZW8nj/au2FVai/95KigSDh3Z/3PtN7Xnjm5Mh5CGoU33YhdTjA5FxVNxCH
ULCkrSxKzgw0ugq5khi2K6DtiY1PueTQlCJpWCtKu+0a+j9FKalPbNpvZnN/GpZJB4kkTSX0jGvz
EBo4UQLeMTBceaZTs8JuV9ldUjuwP+vdHAqHnwKvz7hhCl7XQfSDi6Y49AnwdWhZgSKwn8/yzL2+
UlQ/UuWLc3/S1+SArzw06DlA3mkUD6m17JtRcTWpAaTrQiNKZ3nfTvFreZJlNOssIP1c1ocV7omG
1eAXDLgdjEea/kA64BQ3ghLpOo43kxHbF6XTOnefAbElQ2zPo6inbFUN2f0HLmOmKW8klMT3bo0N
FDxh01031SO8uKMKpW/sUcPJ6LuR+QZ9O4uEHUjMzeQUa+WIN6r4lNSSxntkKgbJ/yjjm/vVzBDN
rK+JGu8xQKt7PCEIvOzxGu2UEaOGuzj4eH+nyl9kZrs1Du2HP1kfcQi5kd0MkbntZ1io/6ka1BRc
vsGNBmVbzE/6uuw+DtNno+XYcl1I2M5n8WbWB1a3sFS0YT3GM3XDYbPUxFUrMmTSrNL/b6XyQts5
qhjiuEYZCFvdCzCBrfRThQJSs3vZ6KTVJA8TwHzliwCJ/wvxdya9jFqtnNnN5anZJv7a879a8QSC
ZgJgk0zo3u8DI/WZ3mTN5LLNXJC++ITMe6ySxlM48iwJNwJ6MweHrT04QbAvpoFcruIC95T9DpUz
gkXqsoXhm6aySDnNIvtr/pXTZGj2r2FO4FMu55PTV1+cdUF0Eakr3q8g20pW3VArtLkLoVvoFyTF
OBr6rjxOy4my6qwi0cmrH7v9Q+7uecYzZym6lmNxGrofCXhBa/Cun/vXIS+diyC4KWgfXtwXSEg7
wNgaTixCgYheiQODyVsLvb4OtCw1InzluZST47kn6ZliL/pa28g4zIVxBDu/XRabZJL/xfzx+OCw
AbAihIkyASNu8tHFUND49QBj707ghhkne3gzLAJ/rm9M+HtOQOL2eClOasuynMk+vunrjnwoofMI
D4ZGM+DXwQC5SvogxVlLPeyRoEa5iteepO8qkXOzM3pbMVxKFQcA7dy+Tlmbu1WoiebjyUW9O+5W
8BmwDcbgpFH4nlX9jTSe99juQ29jPq8BpOSlJBuFOhOn6q+IyntLI5WMkNiv+iSokUdqMg0strP5
FqdRoCISEvfsyBM52nkDwKHRGJXGfNK8Vvg4b85AETnU6tEzOS6ajrnx3TjRW1sEZQvqicnjkeEe
8ZapqcKcE76op1SkuUEZJOll8i+PkP6xXQV0XWep8vRW6hq/EKEIzKVnO30PAJ6dtSX5QbJFP4pr
nL0olIo72Cdo7RCEiuI0WRbCuJP/hjHiKpIhh7HK0k27mLNMCQo/D5pC8IZtkFYctwuNvARMCSs4
8frtGFXbXc+Uo0pIr3kYlzbgq9zYhIooyJ4wTwgsNzh9KvwBAiOe3pBc5b5oqKIUbLE9zbrPI0y+
K1CQLbgWksfFK6ogrfwl9xSAeBa+cO8cNkHL3Q9VaZyGA72BclEmT2oATd44NgcqIXvi9rLd99pT
FuNiN9wIOpB8IT8m6TsAFDPB3V9u8TGKNg4jLFhe3IRj/Q4TEYBU2SdKdIp97wb+NTlWZR5cvpYQ
H6+CWirvcbqhd4oFCXJYZCp1TvAR8WW8lotdH6Z7ElCcXIV+4p6aA0VtTwWjck3CTV0XIxcKhlih
Qf3e+5SGg9En2J6WC6JynWu/LQTSCUW2q4AUkgTUk8VQx9xttVjwxdUddD5h90ZFSA0oHbEsyQYH
yGLgRc2ruSTzVjbnFqfe+3nJhXZnmxC/wuJKb2+LD0w6Mtf2MjTadg0SLfPUrH1r2+7E9UnHrrfn
mH8e2eCL673IwptGbCMjBWLdu+3bQ5uMxb1uyJPmrqnlAbervt4zZB06saJnCPcZ8JZOC9s1vtmi
zrho4Wf0p8lyq8LdzZ4UMnScFrPzp27IPt9aWpxi8tb+AWTgW5HUosG12gU9Ye0IFjOHaFpi7Nx7
nxWu1E1qwWZFPe6pOV0/1i4I91qevSAezGFWus7DmkcppUjHjSA5B12cJcmJpkRJSncsENQAKPc/
RRKAXqFIC/vzakAcxfH8Vq2VAyUpOxmXSTngPYimBXfItNaCcL9ofUbyij+mLtmpN0aI0+/Zl/YO
RiuUnhA1dP8rtxTC2rbMIwUE51SKcrC0G2mZbrwybZAj7gajUiFL20MaNnw4sgDvZhCc4RZ2QLtt
D3ykM5blDiTv16Nb4gL9qzP+0Iq1ZgomATYMbBaloK7P6k8zms6TgveiHT1m/tQMMJPUKdvfhxC3
7mpX4lF6qUB6t9VItUrciJ1sfXFebOQsIojP9OPRrSvn5hzTAZYOJhZsNES6B5MgJzPnUiOpWtwm
AtNGrAHLDIVbo7713Hm9KjceJOnqzudTRNK81ZM23dVNQzDsIiGF+vsrrF6BJM8V4s3OXfP3vDWS
HAsCXufZXq3+tpsWnjTjx3DMMxULZtWC7gAwUggQduvG/FVeHCjUXR8/wN7wBac9G+BPKDYS/JAn
0pORQaVFpUwGnz5UJnbc8BiJrpnzJDwj9vzcRylKS2MqbQP+UBiiQLO7kpqYiLoC49+8vlRlif7H
eH4K/0XnWzPcwHM2UNeIlb+aMRR5wVZSgWMzJROHGjT7l6gEF4qffZ1o0nsY347Wh43Flu8T8dDE
//5qAljS+H0LvOBmFvne7BLvXxnL/gmaNnDBLG3FD69dQ1MmOa4/kfkJZqRqgYBRNyc6NgL5lnhY
Ni2FjcMRE2F3q3cmt0qzZzQX/4OP5vDNf5clTyPu2uf80sxuXGdpXzs5/EIULZ4TRs+4JJTFtF65
n4YIBcOZyBaHTtgO9UydzMPLVWf3rkOJ25wa8HFqkb5b1JUWso6HVMmaWS26YzekRr1hZgsm0u/H
v6lfiiM0VqEP+nD9c7v1RD4YSRg4KuW1mGoMLxn6hJgT01yYs6h31C/OEVDDASlKap2ZLfQsfZXy
/mu0OlKlqkKKn8Zpv18xN8btb9HMp5xYKNKPkCvjgaeEbJVROYW0GA+uQJb6Nar2sW83sNV1CIDJ
bSZcIO/3Yt2zayjGDM3n263fvTbz9FnKrSaYuVcU3CcFsRx9lN+O7gdW523sPsXvkP6FerF+0A4V
qB1OF1FsyKPdb8ArF2qOoei67wNcO1raW0JOvsDv2NqiC+6OrOp+uJVE6saPnUr3r/qnYnrpIZVF
xyjiJkv0BP+hbQu4xXIrPy/KEm/Z+QfLe+vsepgp0RKSlngxKVgUR3+SLAX+91EbNnBh9tGu72ur
4UZkVzGGveJIiBrGg4l44pATEKmj8ScfQ75Xf05CAoGDCO15N8UksZmAhsPLn/uNHF+AZqawB1KO
1+RdMX4snhnL+Hxyj/nKS4e/Cm/7wcsUewhx2MdCJtJGEJqLMwzcfbNFqQEUG1P+uc74jARvwZtU
VPVN23MPIsGwDby8iy2jgAL5B6S2i2UWi2+oiaMPmeScc1E7u3l/YVNGnT5s9YQ7Wn6z0kBWi6jC
vAlxMHI2DZvuRB/Oo73GH8v4zJBnJGvR296VzxpiMDoa4hBgaVgu10yWO55tQrvEiMEe7LztDN48
9yhnhGjZwBUjLbwrQtRitRhGLlTgRfbzrZLmEIkkBMqfrBFgoAamMfTPI0eCK0OAj+wjrlGr1zIn
AdnoCnXXr6Pv4pHMoRxzb0Bm0Y4pQzLvQFYY6H3AWHlYnYazg2eb+g1dfcVrZonn22J8GU6BRKUu
2TLidN2nMlW0NJfua03PRuEiXaRkW5T1tuYgZ893hMLMrm8D0Ofks7mKpXK48gi1LZReNooBReH9
TjU5mU44el8uNW/0Z4YFqqf4f5SAkgoDjHOJokskq0N8oO42Ip7JrXMJxqkbKrMkj01szzVqzba7
QOU3cTbFtIuJB0OjC3hSgJ1BWSMipdAxk0WJy3J/jnog6+thYCAqFomvQ5q+iXaLw4H6EFCu3ONt
uoYB6QrkwTGETql/WATXt2W/fcjMERTNxWt+16VAaWB6OPNFhzNv35rGslkFce7S2wXQ89/UuF6I
Ks8R+jcUkbviNHRgfQ1PhrJUPMoySABk4dpB35AvIOuXLe800CDt6o0Mc7/MnH3jmiy10R7VJNZ7
BpWOxAWQ3lqyBwLiGV19XTzOY7yHbXmXJyZdGRTtp/v1SdR3/5wrhRahgCubB7NVryFP8MKFfiSk
aWeyutbxrxMYenEZTf1IMeSWl+ZbUp9B44fAUVDgxcSu7FYTWY9rL6ZpSJzsOce4SEOeARGQwXdk
lUKU1P5Gr9GG1JkSjy3/hUQoVx+rxvgwtfkf3E6Dgd4TCbqK6mZ7b86q6gsqoWtG+P3txHjA000C
8FYADUww11+62WIAP1oqoRsUOnVZlZTnmNhlYWlmz0KizAH0BE1/543z9tgQXbqofjmNyCpUpTWZ
HokTjfw84iRdhDztUnStXHFiZKyjMRczKN0H9oTQMM6VtjRvdnxkvFjOzVid65dbDEbPjZIN4npW
wMJJOqCMwzrA2+xw1D1ZDhJsTaN912PBZAXrugQe8d8mF6+lIVFDJjFBLgI4csM0BhHdbrWlApCs
kc1b3ysjvYYlr2+xMpuzqZmvRAeDjsXSrHjcaaKujB3Pvcd60tl1SCnMlqqDDiUUHQrY0tDRZ9Zn
kzMbvVZJx2l6+Yy8jr4L3eH6TX+UK3kEPcfHWDG9lZ8/nKsZ3CAnasfxdIuL2Xz521QRlfohOkaH
M978fs1Tb0vbJqZzImKoinKm7WpilJipmd8EiTN8nL7BLq7IYSuw45mBzU0nNjwqEIhgDC+WmR1r
Nv+Ywxz6Cp8lXTb+zYQP5w/ti/Cx8o8FxG/fVPl9MdmLCZiIs+Q8A1pE3B23dpXFU3mj8qkTJTNo
R/RJajYHzi4NOBhOYjeSWQC6hqZlhPpzRjDEOr+cO6G9tPOpQy+2RtM5SEygcaDggj6sZYkbUdjz
MenJXgPh/37Q/NgaWraZMEDSJwU5F0omfBgqGBMDvkUiOxMo0XLiU4EK7wVS8sPjGoUYJ6/N490P
4zb97uEqD2cbpagZffSBfjZnEySUF0PbVFSSvVG+akQTJ6ou6L3FZsdGBBg6LC9cXt1UJRY55XWa
Z95+MJik7KNbDTGd21baPyhQjcvnrvN4SpU0UAzaomHiifkZHnS19Anfjy8/GpCs7Dk6P/UjDnD0
KLMOVLd5yus6Ifk4mEbeKINQubU8uBk1C3+gvC3VS/2PWGgEwpRgXoWyLmLbGz6XqhiimJdgfxVO
PQ+o7PSwcWUj8flfwjAG4QQ+YdZiQ/k3tBJZnk59rxsTuhZosaclb45LtoJE5I2mPw1P9Hv6FYog
dRkQJu8VkdgKd5PUCEIAfI0mLFYCjvhrdpqoet3GIehUx6Ss2VLsTkf/9Zh2So0vYKHuRFz2/Aw7
AAJXaiNsNTBWnsbUYSa+F3W44RdcL0YzagmcbPwQ8LRgYpmTdFj65ApdDjdSBy0wgfLkE49lCp6T
UdYRe+alezAM+aaT4dRgs32a8ourHslOZlF/nJAs8YjrbN1/ONe3SKE3PoTrtH0njoFWNyn1f2Mc
86n2C/XSa2/1Kak6TKa19j6lQh68wVN9QfO5mIewX38inMbMu8RUxRk62zydXrTT+LArXFXIyftC
z3OFLR28w5yCppljVnmy46LkuCPa7KkUtITwSSLi8Zpc3ND/ABUXCZcqprAbt7QWG6u0YEpkRMJB
E5+xiufKN4MEW2HmWpjakj/5+bOuCfZ4F0btjq1Pvw6BqLLDovRUaLy35Ax17UFHiIT0rz9Bed1P
8lZrgny+wmOntxwkCscxwNNLHK/f4xCTpbxWghvTyvBgrZZdnE1st0zVwZIC3DjUcyxbPnyaA3WY
cRIwGJ/9yck3PuFPpoy/CMUG3exJvGWW5PCdMKUSTsb9C0MFmsJsAwNLQCQlENOUxmBQkGArtJK1
rf4upITvpS1QpHVQaGz6J5Ad9oE47bNr90+nSLFHiOzU4foWgtP1rRWqzInjPo6vhUTF19115M/N
CnwmarW8yk76cy0gl+KOMSNz00MWsLh8cf/2VIqK44Kjpgreh41+MOUJv+ZfHRcemOwR0wuw+8DP
QPO9L1HnadFOf6dzO8wYNpCWztq5pQxZf5Wp1xgVcdrpNP6xdux6J1FTaISTJB6SywPeEzuBzINv
Ublh5OTVW96jXGQh7p6rEjSH/34GNRss9P5N+bFgxkNqMJOLIlVkDjXmVF1cGYmzGj2NidGFaT0V
Q4So+2uJltupOFxjtAPHiT9H+eGY7zYE4jU8C4v+nBMmKcBPta2ZH02gKfe0FAW6bUv4m4ln+srF
NXvzVIXRgfcix9SFQtNSeh6D1un32x0lNPJlWtU0EiD3vCKKjydy4Y741pIoL15jef5ieoAe7RfU
2LR1vIzlo6Oi/54QK/uTPViNdHL8etTXRYA/DtS29MF+uHTpdvKUTiudko5o+7ZbL/FoNXmWpChv
MQikHPjP/fHuoM6szp9f9AkYFTdvwF5TIVMssUhGydYJUUeNFkjGwaBgtXYYkNWzv3B0HtEbOTUX
sCT/yI2Fr4Fr14ji6ytM250Y6e3EFBFd2DNSENuMMEI+c5MCCDi5W+SqHqE/DnhGOspYs2ZYLmxt
/921zMUOCeVPsWmcEuQpSMybUVflKuvKe4mXUfZvKZExMLxi4ysVG8OVRpfwHAG4OAOanmS9xnkI
d+ZbvaKruN4OQp0tR67A9hxb8q1gGqfwPqQmhu1FGDz+9Js3QzNkj/kPIu7XWYJUicITXDyAXRIP
xgMKs+z1wgdeW6yczwWM7zTewrkq3mmV4s+WJThdsbm7sb1D63MQ4Gg3dXdg453KAU49ckdG2CUj
BIqHRxikrwVp6EL6P3A854fGmMwlmL2sfJ5qSijrM1oYBehPrMjbtGzeuIPP14NDXX30gS9dwMG5
5R0Yjdiz68AxmJHza/ZQ2Hx/Q+dvigzqMv7Pp/FxwP2jf+evMICtr41xFpuS/pX02vnoLUN3yb5t
rEkUaltVPefaoe1BAQNJojc74AuDr+ZNaRE5kIJ49k5bfCH7WpkOjXCfvj9UzHaGvxltYJ6Q28sA
3xle/cS/orsEatUhYysiUPLy6EP5qFG0DdUNsMrxEJ3c+FPaSvzopduPRtpZ4V+dtTo0CRQLwzuv
wPxDXg6UGWbkhSBuG6LsA5BkznOuKZnacyNwm6dZDY922CMY0SbT4x92sOTpSsVhwMyHAzb4qMYO
oAzsvfGA1tkIY+2DCBaMQeOED8D3VGyfhIEu6t9zaCs1EjcUD51bFHhOzm5rtQdrV7tWCVB5hjWD
zA10S14gjS4fNq1tJ3rWToVNOI5Bk1SoiZzQC7XdGjUOANBAViVRpTGQM0tXBRQzqvKYoiBuAmD0
ilGaZSAQ5r8cpNQW8/E39lLiLtLws0wy+sjj0Pp64ouUXBDsqXA+kpKx1y2iQpDzxJ55L5hqUawY
lOVQSlpjJgivd8na1W0sSvAXBBAiLKTRyUUTkSSYvderTBRcChN6CKIpLm9WXG11GH5McL1vMjSO
4VPiOJbGOhu1AzWfx+5jslf5eCRDQPpm2dFPQAlKsIDIkbRIJU3LdgJ7BIUBdBgjll22v6GUcK1A
JCxUl2rliJeg0e/gQkalzrrxYc9HM0o7GPiGfPQOXtA65kVTa3R6qg67SNWucrmcXStxJqfemCE1
Zrjg0wTZu3+Kw5PMP6lwH34JGumbTQKeU+zyACdrimOicy+pXatTb3bNwgWGYROE0evZtIypslAX
6P1tg6+elHyKOcarTdksHelRghizMqsmc5jGxxRRxXRYcHZJ6gwM5RSqRtM7yDUWi434sA1s84VH
XB6v46SBdPksfoUoNGG4N6IZXT5pXhQTMtn/4GSChIzlc5QkI531XeFDWgQhqlUWawOkPZn54ZLf
KErhKA+FCn3gva40o2/DHgiijSMt0bGMtvY/EWjpT/dNZ+3pHqt6sb/IJc9HuGvcMGQerJ2FAbML
U5IXTbcBiCS4ootyhhm/uBYOBuwPrakgN9bnTyzz1le2UPsvrTlrPuNoUd4sMvOZIR0wr3QdYqCh
HAtzpU9iDZM4IlHKAoBpI7ahQkCxmN/N7iSWa3v6CXivGYTwzNI+Nzg7iaqtRxBi2Yst0tXD7MFt
AwMsmNgBDVaXahxV18dIpuORgj+aJBcG5Nx+X3iCaUFIgpXKPwfNQ7eC02/Xjdvt8afBa3TolzI9
cqsL8F09ksQevWZGMnSwt/F6UrNiZz2C4rRc17UySdR2Pbie0dDh2SqwcCi0nwZhxzEoyiiyQjXp
clVDQ4+E5iqwT9SF6Z5WvMXe4Q7oTVoAafwJfdCnkBPPO0jkVrqUNGVSdGjYMMsS5E9z1J1HybeS
y2VGj0g1apZ6XWv38AQKIsNZ+cjoh4Nco2CUotl7OwxF9OYA/zuwEqAxCxEQSYm3WBFd67qjuWWJ
A3QN2IV8REMa+H/m9NwrZgF/SXvu0YbhtYOtkYjygFYPaNxhC9pguvJyCmiJm33zd9sGqyO3oIbp
ki45L9qb2jLwdpf2QRr74iNFH5ffzqtDJfJuCousnh7zRVRi3yru9xRIJFAhA9+Bl5U7P5Cv1OjZ
vtGqctLk2wgsLZZ/id7HmuZsB2iLEbh70kfViTPfYnqo1ylcIpDuJcx3BxVN//iLqRuha4Kv69hT
axSs5s/XOuWkrfhQ+7qCeC7xoBokumlsQWh4bMrKu8NJXvaGO6Q4KMpB+zKYaDv++1VxBf2eH3la
l4Migf++kaG6Y7ZXs4j9Q/s731626B0lGcn66d0va/2LxsnphVKvGlhqX44GuanZKzBfaRtoh2/U
fKp98+idjQ17cufEtN15xYOFKhDyZucHrLBdazB2M1gaxwTjKeJ8YwslWTOpqXb3Cgo3H0qubSfB
LuDb8x+RkJCde+9D+UUZuyx+15RxpL/YmLwfnoBeDxtURCaO6AXqxrt7TNIgpmKW0hx/UkWED8am
vYtWJpO+oNuTX/scA2lWD7ak74Yu7WEASfcqfzrF9FvG+3kvirqSFbkdFEUx+KUvc3nhwfXjMs8U
6k9S8AQS/t9xf521tkT5bacltbGPQUUXD54GLeXOOM+Jxxkmlzt/KZ4+GBXa0DMY6ItIP7jl3E+7
eY2BppovMR+IZ49JvehQZz9a7dLGKZbONI2GZtqAqdjZOrnYSxCxymzTOZUeMY22wpPWuuOhMUST
H7bAdhFPDhiboPdJGE/yF+DaopCdbbVYZJDIWzjnNc++YN6BZm/c/lRrOeMHOd4xGZ7zXTxVBdIh
deoILHlgt/tVllvn+L66K4S4AdVXaVuLSGYu9y/7xQfSTHy01VWwvVlqQQbkC+f67Esylh2a96ws
qrlFQnmbltLahfDIzcE5TUarILU4CkYaMwlknPcKe+zXMFKGsC/DKXSpgWidnIhuGqcePHpkHzoU
tzDCMoSIVQsFU/S5Wcbr2r6IUY4dNB/VI89a7PN1vgntSvvHcWf88trXqRADVD1vfccfx098GSIv
63m4vAMto4ZunuIfVBnOuA3FjZvuC+4VMMgNAZxwHB1ULo7G5Nfzjp5KDlp8FVRGlvhhjp6C2uMB
qb7G6MhUe1Uu8eClHWk089OTMfwmKzPGN/EwlVV5Gud1Ky4TjbmXOFf+DfPr7rqLce9hkk//mjK1
+/T9JM4zvVCGO6XULvxjULXdzMo/EHFdKCu8DfrN2KC32xTAC0L90R255zCh5fntA7Wxt7wAC6pV
N4RdCh7pZxbawilBwI7ZIpJVrynkWlsaMgNWsgo4dSp7j7KT6jd/qai7MDm6aacgRo6rY2lRCsD8
yMgpOq2MlEPcL0rOrIxrgDXeeYXfUp3kh3yVzzuDlr7tj+TQCLfJlyvwv3YUxABCIpWJ6H4Wi2TT
uLylPaGS6RkvKVEyBrAdPsJOYjwB9BaG38JH+/clk0/9s9PezT65S+RGomvQtk3cfJ17kZlwJLwT
Cb0jV8fKerEVUWmbpzuYiGIK1AUMYI/1wiy7fryVFN7jyoz/1vOwq8QLstK+Zcbg0hZuIZhxlmfU
c/galxWTH1zuZ/hKj1Qv1OIOj2SIB5rrgQ1oJrI95Rmbp/oMYrW+KyqMnWSnreL7Kvmlyvmqgl92
fwF+SzOcfk5ibb09YcrpzjTc6DIDIlTRoiwFBGYV8S49/Y2fk3JnwVagzPSRJ/dDYSwb/l0g+KJK
Qaa/Ar56jTTs4UjPt6Dc9MOGzuZ5h17JV596wBCbfbRRjBoZ9s+UkImzU8PBlA/bNlinZenkJLzH
pu9J3PGQc2DmaOv+xijb6E82dNyDx3sxp6QAO4dQjw1xZvromxklz+kwYf32BXYbIZVxV6Agn6oz
s/VG4i+8JPhnPW1WKSbswnxFMES++Ai3vduISg6rhfLg78rFP/olZHgqjlXiv+IyST99sC1k/yJC
+Pd7AJULieobsOUtDkLQYHEEcTa2ooJ5Prx2K8j5Bid1wR05GfpWD21fZcMXHYrJ7t+Od/X54r/j
MtgHLcUU33FZTTH9PtWxBx8ybZT6zi494uo2kjolG6F/I4KyD/4i/ZS6T31+LU2snZ1tCzkFrPV7
SqCkb1z3gIrs87XGErzEntpHPBgaPx3Wan3B+nt4YTIS400t/dFKgaAhKAb1wd/DpOisjPiYl6wD
ONvIPkKEr59BSQzALhFJ/WQES9964urttphasdsXFwQzi1hshvSgn9XfjxqEjy115dNxFv5tN8o2
+bNmNw7wpwu2m1GxNidN2xlBfGzLqnojimc9kVDKPPZoLZiR61RoLFR/hw2PnGA5Q/kvX2IexiG/
qr8R9eUAkYA4NoeH/Fv6w2ufHMMu52eyGihmEOHqdQrShfU3mSt5hR6/kmT5tZLP56C9ho6PKi32
YiWpodOT7TMsa5AdXlgD/5ut5W6ahNbsbdQR5GHPs3EAzJ/3exGyD1vlfqq34TBnLVey8qoaTGip
ALCRi2cBiSKvTAxkG/8WrmyFjggzi1MnEEM9zMfVlLSaQGpQ6MGuSuM0YqDNDm0PElLCzF1MfmiQ
9gRW+7n6o6F8zeUcUsPuEOwBFegxQzEUgkRHpZ31B2iORjK0aGS+zzbLsiwkqTsBGQRPnG+zRMgt
ZQIbyAws8tsAKDdvtAD3K3B09vW7SZTOOJ4+ILrP+JsWKdPTOt/ReEVLYZOrfs3sOVdOxHORj1db
SjDKWhGw5ZwDpmhlmWfhsQqssAQlJjX56dCs4NuQhrJ5KFjDvpdIF1Ve9yQt6l+opf8G3BgnnJoo
IpRsvlISfZXNRauLOK/M336/TJDDICqdLHAZixbiaHfoQKqZAzncCI4PsYt1MMeL6Q7TGzeA8P2k
tkWKrHy4ejx2Tf4WrsZbporD38BQkAXYCOCoa01Oruz98tNMayKQPANngPsBI/0VRp+7y621YwvF
oh+Vxi9Xm2XzUvVn5675+xxPvJd0LFI5+rLmeBzdvMEcMl4o8vHb56uTTWnKMVuvB090bZxR9Fp6
YJI7Y+78rktSUBWe7ET0VHBB6ynskfJHh6eRPzYqhGeaAXvtiCNn/vJqRSvS8L6xW19tB0HOzZlE
nhgSzgFUpv6qNNJ307eQSxG2ecnuMY/T9aEsT8F7nP1/kqIQi7Bf4nyzf29uQHyaqBpDitfTfeiD
k/P52zD0jC45WId80jl9iDURN+z6QtBjQi7tZhktun2WNGB+/FFh3DJlvSZPMZyXEnbJi+Fh+IfJ
cHLrZ2w72SyMbRtNQ+w4YlsJaM27yd81VaZBQD08O42I4W/jspFfkvRmjxAqQYHXnvrEx5blD8IL
SKwXoTfmoR5uhaK8vzptpXVz007QjPiHmdZXBmgxodN2s875UgMOVlc68UxcW0+6cecvMpcEZNXF
YIXtJsrK+GxnP+MrT3cYHrCWcR8rtzDLUgQRLGV2ZrJoW0u3UkyU8CNRiYBdR5nIWwu+3ZcBtJW6
Al8+TBAuEaARPqA5Wlnay1dJCAngoJzkf+A3jBwCDVJEw3c3psjcffoToQJxd9xbEptYXvpaOssB
Q0mmzlpwT6fJ644ffJtDzHFf7Rv735gCtWskUm/3oHwP6T4b94bPLVyvLWwylqO7Y+xl4pqpSIjW
e6XlGMXDMmAiD8Lxqq2jEUx6T0Njl8bTzD75WxOSwFKOQynoRujqDDYkINp9boaYMKl6wf1Cei/l
hx4ZgqlZp5EM3B9NBZY+FIAHE96D7oVcolutgnt21D2OnhZDLQDWr7cscCVM6ExDY7NVK07TJZCS
gpSuIxW0zruVvKx8FuBD6KNSx60f9rPcsg9cmz81voFcCvfvMnVtYtpH1fdE+c7xublAqfus4oje
p2vIpfFTb4npwau+93wIf/wu0OK154Xe4SLSZwqcPNevOnh4Ik76kQ7UkjFhRVzetgWSvr5pqXSP
I21xg2ZPrr5+LkUIz52rDTXj3Ci3n+PHR0H2UNEKDzftyFBqmxppbfqPLnWzdZwugY/9P06nIfUo
qIpFYLbpd7QQE2Y1gQS+tYovONh4r+WRKSR83uRz7l4ekiEYh/cxSohK/+Ul/qI/pAzSzAzzfkak
CxYQFkIcjMo1i5BgczR36dgeJLW077Gkp11FB66XYYNbLwFpKsQcwy0L0SEGq7IZxyjNpwg7cJMS
KrZiIgwMtr2/C+wshPsZPPhCle7fxeCN1j9x5HLxILDFJ6nIM+f8kFeMe/2EGi68IJCaL7hwSihn
GFyeu1KsuH2UVyIpKCkSn4y3pz8tLM7d31Pkkv4X40+0k1rmw2EVzzTKwlBMIxFYZDRUZF1wrmt8
rAhCbE1CFsKq8bUUp2DFhy0xkvP9QHqCoGEMuJm5XPCtRHSUxZNMTaVq/cdIcKbhHvqqsPD+6fxv
H4a3bAm0sPrYDIeIpioWIb1SZrKnux+NvdI2NV48yUMwzHYTLjkCY3mE4Uj1KUveM2Be9xWdoi+D
rvNTGO1Zy0ip3fbQ4BRK9UQ/xgMs+1zYo6G8KNWN5jkdhzNADyviqEi41U5P+NFK4rhjCYGE16HM
O2d52mYnjvSS1xoQI3ft+GHVyM8aXjB+DrrlEoy6uN6mU+C4ecdTTnypO5lJseMwFwkXEj/J5HPx
RC9934PbKiv3gSemGh0hZ7/Zb5ZP+lO7IW/sMFlLhCegdQVwoJW+Jjeen3/EXXR3B/lacxt20weW
W+rowaMQXF5yQD8LNXPONqhjtJyUqQwQWas5G7RL9gKwT0wg02bOzPfdjbWBW6cZ5YvfN7iwkx5D
oXqys4+OOrLWxr9/C4VGgK31tXtkqiyxTQp5GFqbY9W1oXRlRQQaAzA7hMwTBEkgkVPWNInnQEJQ
G09B8yswcbm5aeo54fWspPSgL5GVyUOvWUnkhj7HMlVVR4ZA1ZAeU1Zqc0KL6P8ouZva6Ndwe1HK
wmm0vTpW+On+gx0yEydKPWoofzVql5ocuWHf6YlsLFexBqEdfdLiWHLnbZ/BEe8ahBI4baTEcJZF
qhbTSEPdkN8YuBq9X2GwcMGUEXUtKIVw89QNtn/A33rzZGVyGIb+anGe7Yt7h7boWlhTtfWvOxlD
gKiE0xHAuBdyMbNf9dv//r0F7M8PFDy/DASdo4NkcBgs/z+Zz67jfP4hHaHo/gXtrYdAMKiOytbo
CMxXwlOMe7jDBs20ds8WOxxd0+wo+Ia2DP1CjX3yCWZf+e9B9G7xsdCqZW824fB8bKbME9YE+3/5
96qHY7pAoy1cdxIl2JBhg610fJ56NjWd+rBT451PqvKSLwLlK1+fpiBEF34ANLWZrov2NOymIFMP
KveS+2a6zdpajQQh9YwgdorOHZcfdHWQXtvzhfD7M+uySgLkPJuY3ZOxyzLzkg0vo+/+w76yuRcW
twYk9dpUc2MT/3gsqu3SBjfn/lOaUkrLNdRTQRHBK+LTrYs3/sGdRYsajN2Uizp8uFVnI35YrB93
SkpGExvGcTFCfHJme6lRy1N35RVrLvjg6ls/RLhjvg1u3vhJQFD4z0hZy8vdZ1yK+yIjQiNHNVGV
QOiMM1hnhiKKWsleOjTwSY5WFXJUMHYU3k2JXyC20UBS4wBgRmUImTj3ex0rAoWx8m5g1cPGKdrU
ixTwE/77V/uGT1TCuHeSGwqBOPbdV8/zobzk4CwMW95dyubsGPm8+arezqiTgnKpR/G6aMSXP1Mh
Bvccru4uHvBhGWZmv+8HsD+bio7aSwJanNWdWJW90FeMpKP5cvfpyVjK3xDHVPi5LN6pgyjwsmo9
4W6VWoQAmxAlvaq1d5ZH6lqJZ7q9gt9mT+ZFM7s+65V1fHA5eN7Motzsqwydoyz5rLD+DawVubVL
Ug30vISXN0wxTdET8FJTlQlalPYYgU5ELQxJMGNKGlHfzy+R986vwvwVm4AyX5xPB8RAmldnvjoG
OPwphgpIKwzbmGHfRedz55LdNOq7aQa1y7s6pkzvSCULdT9esnippgSzl+XrUks5FWQiUrcsJKxR
EULYmOxUH4+uXp+zgMZfXCj0Gj62WKRr/wSx6bil/Uq9xQDXo+l7YvTfiM5LwMcTwLbFw/gF0wOA
hOstUSx/+j5w/6eeT1madoDKZlIM+1DKt4NzM7PC65UNKiSltMgqiZecSj8IVjaVqJBh4deHK7oK
7TIoGD+IbJG3MMJd8Aoh7/pdHASaH9OwhO3A74n9jrTRkO25mkDfd1c2jtFF8cxd9S8NOfdPSqj8
S3HMrhW51PcPuvMDWJf4HnUzg5heo/Gs9H3P0nRplznbaAHjkQoItBWjw9o8GIHSQG0S1Oq3pufs
fKoAJo/ouIuW6hnqmHHeB+bltbY8ox2WRu8uksrDnUL71fHMcvnjaq8lJpJzTrZBCYn3JqFWzXcz
uYvFeAO55a745VVybAzqYAjJLwZOBaSnzSL62Wnb8NyXRfMWe93hiDa79SclNQRdDUA9IkK+NADg
am169ODFd0KMo/xNOHUvQhnJnSpMbodAKWIO9lwop/sIUKweLioXnJEcd6YuDSARPv9y9cK0k93v
vrLos03enxrKoSxRfDabUR9p99kNuYZIvJqpN8d+ecVeIOb46UsSHFJdyuPPGg6l/DvRYzftrAtH
8buYg4vnQI60Psw3yjBE7lUoiHaaXOEyf1ulbm0XOoytfkGBvSFt/uJIX+2aIo8SwW+lnyjmqCUr
iMROwF8+QX9ebcU18BeZfTXpNo4Ij2BKRLLSrmFbj5m2k8cMcKQjDo3VtnmLFXsawaUiMecEm13J
z9g+1Gh42ezKDeKpjxP21asVuGSJTYYc1mAaC14rFmZ3uga/BwizOpZFeTTIVSR3vpprjtH55q83
heJGSefJaM3eBZAxSRkK8A+gt2MtH3nfHYm9ZDAJ0HT0k2ppb2u+F7TvnQ26cbRl0AHC+1F+hUTs
q5Ja5v5LCyzI1H5vfeKShhAuvPh+paxqRr9T8lWTsZoPhIRPJ8oARxOcUhCeAqFk25UhNaGLKtFK
tyZAdqETxoH+5dVo+exGeVWyKOc8gLmcMtpisumQyBU7YgVabm9RT+u5ISs+B25NbkL+bKNEeQLj
6aAAafpQfjkRZWQVD2mYfblz/VALrUk6Kb+deHFNKqdqU4qgoHvxs/UQc2iJhx6tKXahgxrBk/Oy
dVzVuXftOdHtQZRiIBWuLVoh505Nl0zoJcBmOdGsp7BaizXTEpoZPQH1kzoTXUOXJFQxZ8IIChF+
j8rXSNoOCBWC6SkdtGoyG6eHV6FMwyLgthyWmHH8uh6LhqOfw8o361NV17CHmTUelZhN+QTs0IF6
F00nEy5P4MgnD9jrukt7aYktahGagXevPnbCRopxdXpEtNIPMqBPx3OihBGiiSf6pg2wbuN1S+kA
lgSmnhaO9UHoguex/mXYr3Xk2g/aIZz+EE4P/0OFmlxk1gNAmb5X6tnA3yldWuupaZYPHilG25+k
+9xrDDkS3E+Ge5Yp2knN9a6M9cC9TFRGcfuhFJj9soc7jFL5ZausLfZAEyLWMd33SzNnGyCf988G
HjkePUlsb95YUQjzMXABVQCqzfQKTAAiCJibxp7r8cLBtFzhgXO0Z0nbl7UFM0MXzCRMIDWvEKRC
ofyV3l6ExMG/ROqjUiHyMgT+bFctwKJCbEDcvyxamyixg+UcdZZqWehHE5MXkhK9QtC9rR2TsiqB
hpHNnmO3Z+x1/sLVndGv+QntPiSf+vXOjRKIuSxzhHKPnwyoFchDm6VfCb1pgh9k5NnanuzmK+aJ
Frs8iDBdQj5GNVldOaPV16ORfOx+lShAnND3BHDGYVLB+PVHW/XgeaJ3WYwYLQFcB3gm1P+TUZnl
Gr9WYlFXTa2hYlYv3Ew+LWwl3UOsBq1HwniBXFtMiSk2CyzppTj5ds5YRryeRRXZ4ExSR2P9UX+W
KgTyNJnX89KvyUsugbD6addsocLSx+yHGK49N0l75YZbnWIivsR/D3uVBGnR0UX52FEW8/zwms67
4Mujqosq9DZafaVPYGPHFDuRquePlQV5MARsSIauuV9D5vkQxmQy2GOg9nm/OqPQxoLwsQhyuzge
VSRClSXj8DVcF+WdZAHlpwIegSRjj31bITRggNF4vjIxxA6YZ1CW35mbScfBRZoPKDQ+AYfXMWNc
c2qp9BBEDyr6DqLPHb3P7lo7csjM8Pntvxbgp1/iceckFK7E6A40p+7Q6FPE/JnnQL0G5lcA/K5s
IVoAkj34i+34v4s5RQIRnkoCI/h3wskjuiVwDiEKNwA5fEA24ZodxuE6mIn7NYcXzP/qHJUjEZEN
1ibeDIZZKfeqeYmFN9Rz3QEn9zRpE5VKBmLALfz/eNjBSrJVIFu1RwF/hSaBUBWIX2rFFW0hpS0c
SWCFMjvWxn/pI/Oe5+E/mObjb9MgryAJyDeOHHSr6IuqO8OUKXTuUZm8PqkijD3oUq4ZEkG3BQfo
3yWRd3lEWMrVzr7v/mL9xenpNjx/8eF98Y5dUCtPqHvoL7D2+xactQ7be25xD+UfQsMHcYnqqlfq
dp9PgV7C+cOXVQIcifo5JkUhxKtz/2PZT60REU0SMwH27G0MKOq5vc/bWgWfVg5/51kM21+8yVtD
cEc/LAigqob4Py8EaaYHlAJRjeUDYCmbWEUDJk1Jokj0Y7HiSw+l2ZvPT+roAXfqdFEnPne1oXCd
1cmHN6Wfwfv5QKW7e+26p07SZzrb+ZHph74YFhFo9QYoLPvsQVmr6AaFVK24ZXxQCIvF3YrWvrrC
rlDk0sPr/flQNa4sjk3Q4Re/gETjdxWpzWwo1yi9bHXbbfYcfJJAtgH4pVOZGFcMBx3dDXkfEmz9
FqV+mXjJAh69ykwdJ04RtSsHC54YK3vCJd/PFkVk6ZfquQgkcBExD81URtuWWPmgCZG7pMsrN6nk
AKEr9BB3Tuqjkd5UZQeYksQ2/GFO5pIgw+CRpOI8BVL6jvJjI/yaZtF+LaqkkLA7Eth8HYg7PjH8
oOAEvWSeO7UQY5LGaOwb4Nh9IOnAj5VRBdN3tV/bYX8w4aIqBMDtHScDXGm5+BaQEeYRgyipelcd
Sn8eaQJhaIMGHppoX1Ft1Prv65UGrwlTX01VGd4tKdo1Kh0j/Jre98zyuYRlRO77C7HYI2jAZbEk
SwuefcTzBe9M5iezBjocCqlZX/CnO4QZyFRry965rJ9Ub8RxRKgpzKXIxvbutmg8vwIDT/OeiXFZ
mUiDetaDM2A39pEQIH7OqO/myt+PemgL8uDemfNVuxjsR5I2C0u4i3wAsaiozDW5f1kRcOJR18gz
9q4MwSGkoR+YZnrpNp0zI06qnydJrz4Xs0+gJs746kxvr17iK1qdYX4BqhzxmK1FxGl6oZAKvHHz
tFivf+kRK8kIn2iyI9bxqlC58pwmyj/mAFCXa6BYi5gni6rZKA0PqyF/l5Z85SMH3NTd0jkaFrmc
kXLuohEvnNQ0PhDeDH8qWrQeP+5t4DRsyK3E9tJ6N6c8YUK2M4BwGI1eV2Uzc5Ju29B0RC0YHyBU
dlUm5lexrESuZbH1hlouCtSHSjEt3IoPlmfqo+YBXa71w6JJcYaeY+8EPKa7tgdtj12eCehOGvfc
KrSJ8HjcHLKFTpPKZtpnWUUwqEcswgoS0O1jTAbXaJP8iswo9dyB/vESe171p+HrFcKt5/IaTuMq
oRDE5LBLV0EaumpCfGVhMn8TFQcqzN4xuOcZz1mk4z52HYGQb7Qv7r4BpNioy8g3ETQ52drT52et
Fyhvco5HLZpMPEy7MKDPUkJ49cc8M2hWYSWt1jkU+MwaJV4LDOAnLEjoGQKfRMmAzvuUV4Fu2WWb
aD/0c8XEd7dh0gvMSxn3WNIt/ef3qXAmMuE4+vz725I0yMelkzdJpjn/Yn5ykAUKQ3feTrXcOISw
m2/32wCa5ukNMRmMUidQzEENizYly32+tkN0/s4axSRZoNNlNaZnLkh0siXS8YJm9MGiHp2k+dWn
ctnaRIPJfX7n4smXXGw+VpNSfxkdQSIr3+rxxpD771fVYjM4jUg7Yf2DtWADPa/TkpFqHbGz9Dp2
c4GCAR2pDFmlOU2jySwdML361edITwVDr/+IjC5KTUo5mQ8dha8vMVHr1brwuzNP9OuY0X7gR9uM
Xpe6IFtoABI1hKRL+jLIkyNNfbh6O/6MrScL577Ca+vupfYT4IEZUurddwGB9C3lqHPMYweq/ugh
m7ayc0dqk03TDfqmiPeQwZMKq4kmXus+KszULB95aovdPraKFkSLNnjAkdOqdc8bIZe8WwK5ZPpu
y9aSq0chJoR/pug3S1UwHxLamXumT8Yn+p8m5dRLp+w7CFoZeL2Hl8SYib4/9jD6JrDtUhhyUdhg
7xfMCpOer7FMiS2zxQvOxlvnKz5lkQAibdLATZ/jVVZWxWZQYjOrfUUp4jPMpXocL1g/OdJhk3pL
PG9MEU6NT+7HzAwo0Dz1KPgU1a9A7pGm4xcPbwt1zrCdCGTjnO2RPKhWpDCqSMPIO7820+3rPWpW
W18NXm/cb/89/0lRvXKysOVDonJR+6DZpI+k/DRADdnT1ZUerlNedAVua/KeZKXHFvsfTTTXkBMu
kn2XzsWVNaA4+BCvsCYc1qKPqYSd53EjZbeCc3h2pn1FbFNeD/OgaAooCL6Tg5d4S7SlBecHKOzD
VbgwCATciACSLef4j/flA/X56OAKs+IxSSuQo2o85/iG8rRJgfRKSIaPk+zi7BKI9Rvb/YN++mgB
aSITyUPKf8yGKjmi68H2mqO/wGegTGlhMYlDIl2242eJy7YaIRbFdMJDqjsReht1ekILOvTOIGDo
cEQT5hdEDt0xARHWrlTMRkPjAsfvXyjsAbQnimvYZCZ3en3GqaBVI9XbRa2gx2ZCcggPVVPanYjn
LaD1wo+Zgsm54QweHFHPyLKZ7l0mlqXA9OVSIlAbla/dss5UDwh9kdPt2wrepWvZ15sFrVFwtJj7
z/ORXjR2zsIOuW1yv+6kwC8h8cf8zVKO1KMb0NBPct1Hc1XN47Imr4ha/LB3nIdLJz8qOmmWiPL5
gS/JciD3x01oIDWbmUjCzMmlgWkcMmQqQarUR6grv25XVftYe6Z9waIS9/NrRYZ3bBpZ6T/+Iznl
Jx86nUVlO/Szbu8m3FNlW9gJFxOfpTS6j9XXgRnkUvAAH8VIeKPIfL9jlIBzKESjVlwUlEvnngRM
DswI3Te+yNSyozhRdWOTtgbRh//42Dai5OhlEk+ITXfQtYWWhPX8Eu3UXWUd2QUInr6OwyVGt1e4
YUUE85PqmGtd58EJGXsnWtSqIRUltozanTuYYDYlyObor08Bv+UVtF1jT0N/I1Wsj4nJHBx5g0lM
Eqb92b/dDkrZHofQjwrT1avs5yCZtdd4LisXgOGRhM6DaURYbi7x7ku3PsKwp8VQF0uow4ReVjJ/
1YBGKynfqcOB7JEfREWVxaTcTJCPoyvwM6OHrS70V72iV3Kt4XRp5KZFMCnkuq0D4Rgh/JRtN/q9
4b2CoiSrTWjFT1S2HgP41UBM6P4DkFnBOCfs1SLFaiuepYHQjPOhpu2XSbcPBM5ErUr3x1D9rT+f
EyR3EGNosJR5rnDZle/cn1eMx/l5tQcABb/547JixNijhS5xMJ+nU4sjvY4aeHnSuyPsy315/vQu
6lv8s0fu8BY0UEEB4AaYkDSO7QGHN8iBeNG7tPXgPiX4WspCww2ltSewspuV6RGGUsosfCU2D6j0
UIzCTP+MTfUHrTps4wXHGoUXormzRv6lRh1p1ZTsK5maMik20dH0qalaPusDBLfz8RYUcZrEvAm2
PGwe809hIbzSNsXc1zVF2k1vZ6kPSOa3eyhr/EPO4sgnuijMxTDlHA8n3EqHy4XYmfTmgXRYgUJE
xMbwL5D3Lpq/j/yEpNo0O2hxuRnz5ptFcsgmNahTYpNqrvVSAMfT5X4PdhRhV3Xc9O3eLcbR3pb7
FMNMp0k4jQQM2T0gDSYYw3PmZ3zK43Gw1Mll4DHa7/52zbSu0oIK/nOHPax7I2tUjJ5NYc2P2RDv
v9hur+scVy5yg9MkaSiu58ONPmXKPjCyerYskRESIObMcec3tMceyHCHORluxULCD34zuP/NzHb5
DXUTH7JPLn9qcFBJ+Ibfscv2Ry7pd4L+DX28m60EeXgchNljVQxZrz2pzFnlFHbNhoPjaYtWFzU8
poj40nVg/IrcVw4783Hwx5suD5q70aYHZVG8vpnlXn3gZ95i5gFM7ov0/4yipmgcIExrR7wKYFr/
D47rqxX2dkWozgiFXSVo5zQ9ElIF+rtS5y20XlhK5zLMjNXyoeYcjF8EAF/9FFXuXv7U1TMbY2e4
x4WSspS6VdtmoBk3RR5Rl5BfX3t2WRT7kdH69zA+6gsFOt5/dtbjG0OaUWb1+QuEiKn/kcrGmKu6
6UNBj85HJZkTmroUKsiyLx5Q5b9n/4G22dSK9RvJ+C802Zhwoz3vMlGrMKetn1eeNx6zLU2wVLq6
OiSehTQk3bFz2K4MeUidBgsKZ6igFjEa/XcNqiCL0kr2AXV0/KII5UjXy9OfoyQ9nndbhaXEkLrd
DHVCo2Z7JEVZp9PU8FCsGUluA38WAy+5KuP7oW1mG2vIQ4dd53BvSIWpohMX3z40gZlAPMITDSn+
g5plWYfGLtDTTyWhjO6q47A/XY0gERxmm2RoOjMJCFldezvQ1eXtcUX23+kGBuNDTBcCVAsK7pQ7
T+6qYBR1lFKFkQQ0EzXyFqgRxEOd7pbYL8KY7kbZi5ejwlJctsCYhKbO9tOxQv7rXesa0DBKbDkP
YkAsNQtJ1f7Delgc8fcr7+qTDuXTO9t5SWJRY6q67P7bwuQj0Ts6U7KwNAwZ6SNI6008vsflRH1b
wDEGP5PTvMzv5BQe4DLYS27wRVUvybhknJcTmItNmW+TlG9aM67U8wXpF/5PFdbkc5dnyvarw7YF
mBQXmg9dWdUYQa7eCc9y2bSDt529FdtglohPwh7Mhhe3EAjLsmgwYcpIg96tjUAr4hcypRa21LO8
QVMop19pw9k3fpbH4vkdrpWr7n9RhHiQHa9R7c5m7P9rsDveTZQyVcu/jSaIxgohCSF9I0ufM/RL
q2e7qAoTgXRlekm5n+wVtMtOW4wXyf5z8o6N47AQn8yVbvORaYsXNhpaFBaIFlRmBvsPSTwuBdVH
HN4GVy+9Tl9Q9YycrSQtl+YDiscK2SKP5VK6UV4oy2V5IqJeB/jRGuFC+h3JmVaRsUtjXG8C6yBE
LIk9WOdzvM4riQ8ziJVz6KGKIVcXoe1/xyc2eEeDLTLNWh+13XhxceE6Isz0BIlkbStdFQjhzEDM
Ji10rfcPnlYZ4Dqq8SQlCM9Cy72OhILlnZF3NgZhnX7KYM+J2xSEu2itGafwbKyr27JOfe7UfYjb
s2c5LOIfDqrbgRVDeER1sGmN3OiWyAJrfizqGcGNxom9BUkuK/GgGj50eTLdU18QcfyWo1NhFth1
zCIjH9SvnFIjBQZkxiztS0pZekq0hZCuohkkmQyBwBeU0l86qfwjt4X6XtmR4anZWlBSDElne0FV
SR1VlGCHwJXs0ZBiR+F1OBj0xDlDcCWe5nlaartFFZPpIijEX1Mwkr4Ccnwkx5rjm9zV4SSsM/yG
7Snn6WJw2/eMXclPSO8oZ5szXBQBOgUAMzjny+ioTwPmT/dlPH85VutXrIGX1lf0j9M4m6meRfdx
2HQSua+cMOAkJyhRU8g3+VeddHFQMq/q9k2LhfVD1+7FeBxjwZx7cQWDO3I5Or0GV58zyRwTd69F
9Yvz65wp2F2Z8MdTgANDfp1NsRYMHxyDjotJQ+Fw73PGiE//yRgXnCxCq4r01YUZHVAXn6tgjH8v
rMKphXOGLZPHdO/9RW7VhbzbnEVLfBc+OinK0j2WbgIWvFCfDGelcYYBIV6ZdWg0Zf4blZGEWLa3
PyxYUsbtMu6EOgwtPJbZZLwi5BqdY+HsmIUMMbTPfeLWF/i6UOvSblZNT3c/CLvGPIkXnBc9EHdM
HDdYmXP4Y1UGPhYF/5Zb7RjL8osKVk8fr101bKr0oa+zM3IWkBS4s/G3cJWDEicsTCj2m73LYutK
roU6SDJ72t0UYuAQRCd6PVp8P8pmzBJiLdSgXKCaUHlPgQP58jVuOv2l/P50oXe6l99bv4zJf3Tb
BBUlkSmVKSZjPsQsKwQHiHOsJ9W3GxKwKjWJtTYzyvCrZH56LX8t9rfCzyfDtsGPcgmf1tkAGu5/
g+sJFqmjlV+tdySQYH/yVAsClhklJUMcOUNK9q7UdTBotP367gjU9KbYhmTo/WHwqbvN/n9IIZe6
crqa+c8ctbYcPy0ws1o0qloK3ygmHMyad2AzzmIxF2WPpYVhwPqwFxvx6RMAGOQzathpqZm+njGo
Q9mEGwkx9uilhqxgqU2SLAAuFXjhfmMOny6KBZGchWlhB9K8ezTJ/iDG5F3UeDOGS1Cbe0J8rKJH
IPXC8/hDHO6NNOP6e/ajAlKLgL+/08tvDFyYX/n9yo6iJhmWfyo/bTaDoIn8hf+NBHEcPZ9EjP3z
bdP9oN2u9VWPbyKJnVz45bhy07mF6NyHg7KCmuz6vVaLGxiwgaLgt57h48oR4a2T19vyGKCmo9Xj
beJqlqjRHLKAjKQKFV/KOYvxzzpxUQfHIsV85hf/zcP8JAi6yUHgOFl96bkKJNyIil51O6C0bdY4
BnlTxQ5vq8Ix0ojRHivqMqTSmUMl5JM6LjR5U2enjJlCuEcIRmkWUIGNodVQ5jVlxv0M3QHXDWBS
nvuUnfDzFHN2una9s0pGgYHTmfGtFWzLC85xShgMiYq/LZo4wKdd1N47cIndH9fbqky0WySRRw9O
UVi47A5HpiRgYXv3rPSXdAT/dgrLJDTSJagmLB4rUKNf1RsPKIa/cuknGb6xXkL10kuBF61QN3si
YGONH4YW7+ynB/pOZl8lX4p3I7qs/iMH6YUkMnvHoHG9MsRwXdJMON/0rtzZ8JUkagOZgrHHweNk
et5tqPKL+/kzGcSR0dwDZQ2mUnklGw0WWqJWUfppb4RiGEQ9Cioug0p3NLoiDZYv5wDkoKSQ8YVZ
JPjyDIn2iQZbO/TxLQjgI1Vc9nsklbOW7o2GeKbOH5cckQZ43oPIv51QRdCoVae5lpeDsRfAIN7c
GP9wrhX+DxtJuf0ZrKNQDem5kw1FtHMKR1nFFJAo2WxwNYI+T5hW1/3h2bhHAa9cp7wrO4lXM8TG
j+ggpsHYrHqhaJY7egm8Xkh995aKZNy1ARMNSQhyFUKITRdkdSoskKKCF/5xnx4GVDgH3U1jmJy2
NpoF7qV4NGvjUAOm8VI2qLtviwdPLZMUbi1WR28yTh+fFw2dAfSSFXvKYu7B0MvLwHA+tmMfpS8U
IbdPvva51xK1fYcpHSZrX9OubJ2MymZ9GKoQP6tFF8NhKnI0U+ZRjS5J2q2Wpn6J6YZ2ktAHxLhj
NpaOfodTEqe4wneorJnOMzOb6sUc6y4m+nsYkf5mfCKOHF00CPRVeS3bnvOtwTw3aoEMYz2c1/ZL
+wTH93saZeiSw4CtLXhAHS+yXSe1tEh6UTVgi7IGwi56DZEKde0YrpNEunycGRYuzWU0DARJKmJH
9SYg8TTUH1v2icGlimUipMB717f0gcwDOiGSD0ecWscVDGAbcc5zfRN8eeMGhimQUEYoraQyUnoY
1GRje8rhHA/fAVqPz3O36OwiNfc0AoUjZ1l+4z62c3Tkdr922nTutm5gV4nwDikAWkWGhRxVFHQ7
5aDiPOKqFw9luSgjIPjx3iOxzbJKdjStFdJBolNOwWpPzwCDt7f5OU9tbXzUg3ynJTt0WpkgPzTo
EXMJ16bvsdwvRLAXnA7ffFUmE67h47/AzRhP9IWLyv99Px1lLoQWbLCalCnkB8QCcb2LnaEe3krj
YpbVRoxfQSSlVPCmc8mgFnTsEQyS1i5Fei3t24CUoR9zZVAYew8exfzrbZVOjHfzJti18mQ0hfPJ
aKfTps2SuL72UXkhlTcrxt6KETdTUPg9dzDg22t3wLIY6cbBLe94i3V64n+Luwtb2W9bhLfootxk
3XAmNVQ9Eok7EnkwObrwACRFKYIPaQqRxsJvdk4329+naDGgCMGdUZS24tIxvBzaRFRfVAZ4OSdZ
tMzp/P9oRAuzgLOQWeNjbDBazu1DWXxINnjOEolS/et71t4/x3Ng8HbKMjmAeLmq8fz4Blf3MIQI
bi+rWiSHcLC7wrFrox4DQbUECZFRTxdyPxdWMeGKcnAszTnKY61qNnB+1tY/4qsz4Q2//XcwgDVc
5Ln/spTYD8QWe9UzWXHxStC2E+/vW8X1Emimm42LjTTWFr+nmQ52F4gKbxeprA0l/od1ak0b63lZ
gtojPwmrDvu5i5exvKNyLhBk5cFyNzEwrPNsTLsL4ZORUVdBeGWiHkcebGyKl67jESuweuqCpd1A
kjMZ9y9jNeyYDUc8dlTFsc5rhbAQLn+oSbZGfwVqOSFvn6EPRogUYKN13mk2CPvqKdHG09Ocbuae
X4Ns7WVhPSj8CBhZSZ6PIXnUeUA1XrRzdyEysPWbHFfbZ6rsGHRgZx8Pn0rFqkwtlWnA98Fke51z
oqj0w3GON2Ll/FAZkgdRkPuC6rO3EM4dyv5zyRZSI7RdIKXtEAPgPRctK03CB4toN1Dgj7jsmZrv
8nATrnWMbliYXzOJvYh7Eb3PZr8EO0HAbMfGGoyh8kvOmnf/pQLytycIX00EVliPvfoq9o+bzMf5
qCUxulZbMpuaS8A232L3T6qTZ8zOowIvluqZj4ToBiSzLU9amScbTH80RivRQWEdMsdFubY3SrY/
RGvwmOK6ZtYYpvx2ajKUFZi1ceD2RP4LCqqp5nuSJjdAicMDpYh8adkYEAWRzJ6CRZyR9JmpkD7Y
D9Z+xRb5N6M8TwLAzHxRqVzH3I11NLFpkaaM3fPJfY6vlXCYLZRXsqvu4Dir8LxGq/vB2W5Va4gr
Vw22xcLCJYEVr2fCrmCyhsOtQheitGjiZgjDnenlqUQQkrFe2Zr92FEA/iBFIOkN4g9KydBvTwZz
XetcqDs8RaCbpgC5Sr9fuJ2nVwwt+FPUqO4JdRB9z4NfI8hOt3fS5DZTHkrYr6wmASnWB/sfzDGr
CFvHVNR6JPy0MlrjwwyyKI8TrxGbQ41egKuWWqPxo+Xt8JVTP+f/zeJm+twpim8OpIwshDcjL3at
0TGlePplbpgr92MH0wCHbd5T86g4Bh3+aZYSvesXFcvvi0ifOWuEFLRJqNp8GOu3ewNzEOq85Ncd
Iel7nlrJQX8pcwLo/5MzW5o+X2+EPfhjQSmwrSIKiaa2lqR0paN4s1LdHRv6/MODI5bHjZH8URZm
XLmB/zjJJ/lQNzBfxaSzOiHm7rvtyPK5bVDeU0MD/ZQSnEQofIW8vYgOEIQZizFx2DguxSALu86u
RJ/FvBfR5eh9yrtCD2PenjaN1kWeAjntzhx/7zaXARHXbH+ihgMnb6anGzOY88Cw531haU9JVEnJ
tRwd0gIDsKuMvhy7ozmQioQW6tXlSz19IP09TkPPZFC3+4yq8WkkdqyzmmSi/yTGPY5EdtvzhRbq
pLWb6wlvccHkES7XJagalrRm15vweJzBQL7hOVxa3+6ntx11eHrxxoFeMLUGxacEWfBT7iHO6nf3
EkN2+Cr1hoHP6ZqKApqvaUo84PEsXsNg7UYtjia+9CTjBsOTvmKj43o6bipP9PPL1i3WtFR49ZoF
icgSZtrR7deDLs+i9Yf/5FOs0Aadqe1ccYFP2FxBRJuSAQgf16T0H6bo950f7qIElKsxGYbEyI0a
nPdqL5Qbe5mHklCYoZlcpfF2dShhLocUegW5eEBhHAReuHknIJ/aXi3DA8l7NrkLy++qwiB4sbcj
2fO7CdalurSCkFTLZK/CdXEghw7XBIDouEKEPeJT0UM813QGRESaIWWA8aqyUZVf+sgoaWNvxxQz
dAAftRzV7rSulz7XWtm4myVsMGxPBavkWW44pEnwbQhycZSDnKQ9flgnU8Y7H0mxQAa4iLk/2qb7
dHIywIBc51f5joDiidH2WissuH8HMs0vFwrxgUcf4v1aO7DHxJ9lKyf52Mi/vkGO8H8f3w7t/hxM
IjGG5ZAhfZtFZ+OJ77cphpQ2haPhtTtvd4c/jLk4nFc3VwhJ+fCRkQ0GuL+F2B7+PmD5Xy+10ti+
J/tJtATcJmBq+EeVwmfEn/izrTD8JztQYHHmdMKYTkFHy4EtD4sAIu0gprkglmkpwgqyAWCEScuH
Pix3yGgMxMA+s+nzrmFu93kQyDDBmM46+tg2otK5GOa7eXbL25DxRhaNeWHYiUzVc1/D5Gx13BNo
RLqMZmaDv6qzJSo3HzQzzQAZ+uhN1pTkLtZIPghe4F8IqhcbkDIwi+5JDYHLHzfLRQAemtrKDbCt
PoqCdx3XxfgNbl/+qG/y93TT4QXeL6V+sxN8eIimpp2GjJjePp23NuAUk1NEM+H9xc/vEKylha52
kSxLHvmPDXamHfT33AYHT8NJam3iI4OmjPX00TenNB75LXFfRQ9RQWZ8DgnQItMjnbaMf4jhuSH1
JqmHQCE1RCZd6afZ0jbRA0gLXB4tgcZdtmI4BdoqJbZ+vwbj64tWPDI5vKUs5NNuKiLOoHgp8xq8
k7uSnydPrRvkuJzUG1uZotOSt96BqHi8eOCL3sfb3EcJydo6U81eiOEgYpmftRZN/ecPqPu8xn6F
Nt7qPyjp+w16q8zbyAmGkcU8yspGatua+HsaYYY6ioJmGbkEPTVAYXBt8wLVIE3v6TKT/piZPQkS
1WUY9TfOZR2mWooi3yeCKjQk6vS1qjPrnSSqIFTFje4ZpK8E7MchetmShJT9SvEDMmCLE3s6f9wp
G4lb4nfXc45PMkJlBqvLuMQcZOTpnJ5zjLelx2UdKuRk4AohOQEu95BhP/cm6Q+qTcmXWS0MMDi9
BqPy7cT0DUcmf2kqx826USHVL4+9wLXPEdPb7M19WHcCW+5ngAZ+O4y2dUZCOy0T2IRPPmBq2ABj
xpWYdX4OGKZFRKHXVXwbsGf03qqaN8rLeGKW4fHiWZt6Tvu3sEfhtzYlNs7tqszax3f7emc4dFgH
rV+GfWLTxw3vy5y2od1+MZEPqtdCO3mFKT6WjjmNOWx5nHHPSzZuV9fX3h4/iuMuY4U49p8obTSB
4Ko9I+rszpYZPUjs8tzMKrUwsZ5c9A73T5iVzzyBop/zkHpwEvacseYfkyOoV8DeQBEYsF8SSfQs
OMzspJRKzx4p020+AvuWfSW6AwIrtq+Jv3wyrGfUwROpiTos+tKD4ukcxfD2gTv6utHN2+S79Taf
eEBJs9oGYUWN/LI+bZdLQv4IcQejBc/895UsDRFmVTNDMNYfFWz6IAIGukQczOXAINz52HHDk9kU
2ODXcQ2Y2x2UUnPqy9Ut3D2ST0eck5Pp/H87jMao6IyHg5/rdm61ldy1/eTTU5NoJdFUFY4bS8IT
JH9YOTgZ9YdgV5xGEDKR4j+JXeuxET6GJIY7gSxI7xl6gSclDHvDqU6/A/pVOs7hGMmsaQf6qMCD
cckJIgvtrAEXrUx85CTb8g5QCMaN6oSmRzPlMcK61QdJdLvxGcp9oRyREhlcVkrefxWZA2pa7ABk
l8liB1V1XMCH6ngkpUYWrfdMGcJ7dfYCTBNevef3s8QmrIyVpm3ENU3sT0auAQW1Bu9xHQhnoFko
sNTs2hCCOgOTEMpGNSQwp/U/WGnKTZutHuNWeqV4tGSntp2Omxm/n24seUOUc9iy6dzbaU3IE2k+
Fz45HZQOiC+5PWmhej6TeiX4gXjoOnLeoe4Sq3bGPylRbVCwdTtQiCKR+SjwFcRDHan5777m1a2F
dvQTkrdJsZ5vhpw3eTRwD4+c4HFetvMyRtVg/ayTL9EHzIo1I6QwtzHBkVBXjjyZ71PPpTMH1eZM
7yVjcsx2ANJ5Ha1qb9DYpokU1a/Ze1+X7iGCa6nBgjFMpVcqxUbof9CV4iFSIv8KXvhAMETGehK1
P3Q6oz0ZS/nEvcrAPoz0mb3KhxwJPbXKjnNOyEb+q+LsZ0Nj2mkAE8/iqIFjdc7bSa4qbM2dpgMN
EmV1wkS/eSGkUT3zk7Scb01x41au67RvTE0jRiWZizYOJqIb+TKLoSK331m61+uYoZ6IZA06Z3nc
jihKYP+QpwvmjwVa7ikbQS10uGeF7TebUBRb4gLN10iOv/weNWdPrajbch8IEIpyJi7BuH34x3wg
ZSIgy5D2OlTCd3SUrtgfmxk+7GiTrxl1gkypVOMEgYFi688mLH486INlQUi3+sAx5lGzIrJOvRn3
rIOnNhXV4/0wD72pKoMa+p1DBHvGhj/+4nkaB8MlUNuc6aGkX+d/H3aZfQckrx2BM5TOSUFqjFFe
dnqVFBp51Rrd2iwdHt6L2Q9DFVOfBGZUpw7Fjy8egKKFmuGbRqy8Pp/NWftsgFWlJRhjHlltV9JZ
6uChEr/BdwQkRKk50ht/dC7yAAxnOWBmgxUSXutGo/4EpGNv+2L/LuHxngqT2xO0JsUgzkfZcMMi
bsm4DO9CAuBsc5TPbgk5HDk+c+cNxNbZKXszXlgLP0kemxf1Ac9UP88kPHWDiZELVNiZAN8JTUcB
UgMyHTAzF239QYK3mTAlmnTy/uZdH0LesaUe8LPoUE2s2P5iUMJbl2mY+lUjZphmIBP0QFEK57ph
zHVHxPezXTJkbznoFvMw90A4DOp+ERKuV/2R19+qTBnuqFxJFHPQw7WMgJgpdzgIij0hRYkYED+o
qyyBJKNxd6jmlDhTq6w3Z9P7yxwmacCsUwXgIbxCVIecMk6n1AfudidPd3o7GYfbmuM9oLI5YTUA
9Lo47W/9GEOAoQcwcQXSRGsOnMoDFPzaxNkEO1rXueFKllr9iASDYZJMCwTtWNkuz9Vdq0Kwm3xk
IkT8S3oZy8n6C2NDOXz3Lkmz6y1YukiEeuqc80Ktk94bSY/EA8JV3vA0N4RPkACinh2y+f63FsJG
TpIF1r5XZZXDVnVbkqYLZMNqzuxOX4L46s9/hQQLB1AjqNMdpRlf36zUmgwcj9DbxOCVthXZlIwW
wEnlOBVHBUWla2ybkEtMHf8fGV8oYAiaN1EbPyDsRZAqZ1L/0XVwhGx1FBjA7JtjyxQIp+9FulCM
0ZqM+o3ohzY2m414M/zIMnolcc5I4i4MGb3Yw0ffUr3/KWt5lJUeGeK3fv57nQMIXoQ+EhiwMOw3
Lt5CQBBupBuUoBqm85goKJjWYkHAURmRIJ8tRhAEaIBIwPwkFP9GDRIujHQDCyqMF2ySiceBU7a+
pZvEF+9GVoeDUW5mp7iQ7vun40UMtv/wHUVJXFxlxW0OG8lds1kZBBzZQvT7ZCDu8qbPanqhH0d/
jHgznF2Bpe594HEku8ssuF90os83aTbcYAVOseMVvCxTiXwHU9syQzMaRJvd2QNzKlVBXvCwzzRk
osNNxhq46/NfhjXCkOlxkgr0m+ow+Xl/9VlN89SrYSqKI6sj/rhYpufHo5nB1YL7WRCMOkF9Hm02
1qHisKud/hJanKNrwBlAIN9e7tZXg8T6R1ggksA0ITqeAVY2Pk0TBqZ8n9FIyriRgPGozGtXNDfJ
y+zZH0yuxcML2YhWNbnjXFuKdLzbYq7D5/eOX3lxxN49Uf/NtmpPNjHg0ZpMAaGhtvao/up3hZdP
zmAbRrcP+V4ZWNlsOJcDud+EYWYPQNiCsFoK6YzHw6AO9D0hyfyO8VB5RcQxkXcOF4zSo1lwQgZJ
MX1IebZEFciXP2yfLwDtlmQYIDspZ03uzdK+2V2vZ1C/ZoyT/Vl8A5ZCSuBAd5uVTaEWBDm1+EDQ
rs8kEAa5GGCcp0+yPM145iAuzzxfHCKTvvzNy4JiEcPEhTh6OMsyci6vaBabh0oNq1yTFH/FTYL2
DEW1eC+PpbQKuENk5oaibMpUtdSnDb3E6R+nfsZlez2FlzmBfBY+0+WnzqXzArqje0j9jItBPMtw
ybZ+R//BD49syt05DFOJuDGn8ExdBBhJOFEVQ7NqwIEJJdaQQkcSr6OErM2XslCgTT7MgwuJr6pU
vAZbhu6sKTAwcwv5t4WPrapnYG6JUzxCQXlS55PRSFIy3IjGCjQL2F2k9AextmvXx3ESBEhY/988
uhmampPzkerf7B9ZUnvRriJq2qkNfHe7m5LK9NwSeG0MONVTW0EAZdn+0mcwOccnqHLdQyBvBFTn
aSrN6FtfExYDmrDGRC03ykZNNBML+ukiTwtVkCEPOFFCbNhHUy0gcGUMNC8BdKSTpSwvFtKGOCfJ
g0TDLv6Duh+wfVRGnP43gnmDtPNlq1VL7KvHatERmSbfR3HkHnVgtQ0CZ4+9oCE1LfjRTXBj96U6
U9k5BfiiFS6c7trYWywKaSSi2oAY0QwIb/WgzZxRAfkigNxLnJhXkg+KOpfXKqKlfgX87Uhh7GtT
Bz3gvskcnTNxbUL5U19b9ikNonxpWEujci3fURsCjBwhSw7ttCZPjg8CiihKhKxDYV7tYfu+nMhQ
9cCyIHBTX5+CF4mJ5+3jbDkqtzg7F1miXCdJVwsqqjFceNeuS5KF7nWahDt+2hbLgbCtXZw0KWuV
PiD5PJZ5p+ZvPNg+zoQoZYDZ3d2HFjlJaks7dsxcTn8evxYMDBZii3crK049rIw0pBTSvRB99Krd
wwLo3QLW/6gmyp3RYdSeVD0CZbaCE5zdv++egNAd8uSOqPUUxiBVWDjJtPU12YBskIxcSc5aQS5n
N8qY7ek3YByqbzWZ58Enz0eQGS1RI2GLPp67bYYaPzOT5SMOLARDS2CUv0PGRAR8rWoMOlcpMaNz
WOyfUGNXTEGskBXehG6sO1d3ikoRanwcGgamqk4qtDRcVwF8p6dTeppH31x9AUC79YADGbsWVCIQ
JiXr1rxwBbmyQq6IU7ZtjddJqhD1DEbM1LWbcgHPd/GMjlAeAPYZdbxHzQ3zEBUYSdVoD0fCR4KP
SdEoel7T1b2AFDh/UslmQ5RD5ZLIgGvHcO7ZFrgoVeB1tjxLVkM85cxirx4JYYIRR4bGOpIBusFP
93WPiNez1krWrp4tgASRL0SRJRuqPUPLuazJfF+2vj//CwdJz/J9UjFehBD1nKrEqkFoVqKNjERj
2puBCcMnRdEBoRKfO/Eino/ZzONgy6oROPHckhQ+bbmZzveL37ko5lJHOCFNJrbVfdU+qJXRGtTB
2nbySmqvcfIhuOCu8XNpWmosVBSDEbcdXp7yCzqTy0Sa7gQ/zo2DIk52BF3zBtC2PWrr7dOUcw6O
jhBBS1+Ddhrj7f06hKEhF+EME5KtLS5FNqffsf6TPIKVAoPGSRgI3u2MMleTknEz5gBuHFO1g2e9
FUVCZH/mTYF3y/nJTTDBXsvPlMnZw/iWmR59OiNDMRGLYKPGGfT/ew0/i3+17+PBVeDRUqObI0ga
dUP6aTyK2rxyScFKGPJqioQHj7DpAH3GTr5E+YJ7TF752oF/RYz/+MSD6+Zl6EguDXlv/CSuvqmh
UBJdmtfNuEjDZF4UkOAVR/gUYEbZr8cTbdHMz3flAapjkjwhjiYrEXk8Cr2ieg10ln0GzXfw02Oe
yIzxK2fswc0BZ+Z0oW7VCI2R+4uS0D/7/lFGhQiffEt6GTrOpTmOXkDQOVgC7RnoVGw+y54pxzcp
tcq5V/ssVOPO39VSCB/GKhQ9WdDqe8a6NY6Y+mwwDTZYdgNgJ/nR5CuS5LORKMqQwDmdt3Kg5M/i
wqZi46AckMzIrqm5wcjWADD22QlO2w8vnSAMpfr4FtgNxr/HHUyYPjv5nx3bsQfz/r5vkTSIu45M
7RD1vK+WcTNFUK3mTAMpfsEWeqG+7ke76w+8LYKFDo1nAl3w/mXPeeaR14m1Tiwp5L5Qj0pX9hHV
h5MCYxkMeyKB+rvEa3ePabo7vbbmJa8ry0Lqymt/EHChxNIQc0bMqh9qXE9IzB1UxP53YztXpATw
0nl6XbkljxAazuoVnKtk5QEQvKxqnENNYRgsYEO7rYL/KHJEse43ewfw+u+pDxlHst41FD2xVoYT
aSU2AJiiWyciHnF47dAfQoWO2ZWyMc3fawm5YAHfsXt9KT0WcBHrI90D8OBJt9Yw4hLPfhOiRW7i
elaHY3J82yWhn4yDk1HxwkN4k0S3howQdjG+gGkC7xSAABWI575u2ggPzRyELgA9WE96ILtieJ69
bdwZwEZYGCZ+jwl+1jEw8fWtNxx4qcqcCKnjgodRqBoNP/tgVA8HsrrAeMRGwWMDOL74YGgXsn79
NxouGMjb1cqGRgEPrZKyUSS1mZfxsQcz1bqCIztS0dgYyRbEV7Uqh0xtPqJU/n8t353VCyR112Wo
ZUrWCK42Qkfv2w/P2U52w+WbRCVpXyYxQfGTDKBYPl3Hzwsg+zdG4MxN08mgsvGPI/nwqCbw6quc
jn8/KdUe36aqmP5A6of2ZaG5+lh+XKIMA8sjO7OA3x0q+tJAaEQCAJBjXdWgsTYi/FpDe9DDJeZb
0uv49yp9q77hmdHfx3McUIfPCHR9il8MSwdIwWfNADDdARLVskDJa6lc8AO2t3sG8kVheLSJREZ4
8bSVmSkKmLZCpYLnNM4RMmXuGoRJzybcEfwMliImp76sBRp5EvOf5WG6Pv+u0As+rh9wuw/Ukrsl
teOLBSWSi+qXShPRBLARN44EAYi5abXks7v+Y51c/IWOsANEIuro5sn6hjOCfRbgzk3P0OFd/MPI
e9At2ifUN4nNUvLleCnxNz1nRrXY0e4Xbg+jZRFEIde/iAi/wzwrswi5A2nk81KFAwEtMPvKdln2
5lb+cpMfUMeWFRteSk/3GkUt+on7pa2r0qBeZXcj1D6zi7M2y79LIDWmgiyDJQW4x0DKq6RQ4Hy1
09fqehpNglXAwFB85sSX8ou1xizlvMDbJGZ01IEGM7qd68YPLVcMoNzV/i92G6E69fcNkfjop9zY
ce5PJ0Orcuo702JPK9XmYynyXD3eW3DlBoV5YAcYDINNy9RAhLkzbzM0NJP14v8d9avei3H6Xjnt
92aKQge6JZSMyNmHafTuLusLSoVQQg1lqnTANM7KpAQxs3X8coibMEfVN8+ydz+1Mlf9q80RRCUr
tSQ6FSqqwQ8wD9PWA6iZD8ApF28rPfQlh4pUieuySGKQHo1t0ahrczW/82Xy2TVubg23Acl0FFIn
0SLwn8fcPqtefTXR1OeLYCCizaEMxCICt1BUuvodAsj5fXLoaqGoc1pVieFlAnpTmuRaQ397Kg7i
ryBAj70MxPm2xuUS3Nemlpaht8yjexrYbE/4+r6lVky3MtmWVR12QwcWjq5xpEQ0pMOsunxhZ/jw
/7jAx54EyDtrl2h/EqWH1CFiU1mn054ByODnPA99gdflu5cGaI/sSHKzDkz0E8XkLY4fp3xbzqgT
Rbe8e5Y2qJze/uRvRoEw7QOb9HjOlqF46sBSCOZ49ZZ06/7+wkhQfVKgCRjKqjnS5UR6NM87Cn5M
oKmgvA/2rB1/jFyJrRNy487ACsXr1PuhgxiOuI9BgHLf9HEsddmhtJUohzbpR+shUZEWnSyx+F/w
SzRWvnToz7B+8Yvo9d4Jo5NbFYeF1mQsWN9tNiW8HLU8ORJEAaIXQddd4Li2jDBVvDjGzt5AlbzJ
2Qv0vANuR/h0MfF0Z0Vp/jCa5bjNEJeMkeBzBqQ5ypwYbHh6jinxjzMdcvN6CdUk8j3BG50pG5sn
RG5DolQPXYy1PT1gvGAcoLypU2EPWK3/1rWZI4NTZMZcPBZXkuFqzFSo/sGwSXJ9COLZq+sVP5Pi
Jw+nJLqv5bpK9GpwJHI15XK75PPkeBFLFvWtAA9GUKwmmV10ztTxAFz26rNVd57Dcwur+kMKpqHx
S0FTIuxhhFBsFi22YUCM/GyeCify7cD+DcDar+9ZnG/bHyW1WyGGjqlhEK43diqIcGijD7rn6xy6
3pLGMrhtcZeh3q6r465TAgegFFLrdxpP2QFp3W11HKPAFJkE98UaQX3Soltx/uBl03gHxFMa74Oa
icPaUpYue6EzGAma35MyzXLVBhp60/0ML9EtCs5hbOUA/FSRCVF76elOUFhEXiV4yIvd/KzoG7bd
O4TPdLjeNyUgKvy1yUE652Qzh4d8Ir/lW8PJXLMN2Ez1o3kTp6uewGgcNWQz5Uj0nlTt8DSCDpPE
JVoEaEiZUU/vwLwZUA9MDZbdZW8XL6norpsfBUHfKIpemI5K6xizuCNXQzuThGIYIwCoWfyreqhl
rPTeuUoXKBftuesvPBtsERPOdR/COL9nOJvbJhdLrOSKpFhD41DCTsQ72LyE7VIZdG4vpmNAe9DU
fiY3hNiMiNSPHui9nb2LgAGHDGthA39r9BW6XVW5yrojA92tL+NFGmeLDh11W6ELYhq/cwygpAvv
6AyhgUpvECqPWePS0ivEobkl0KgdDEGK21f9jF4CkYr4hiirPosM+J8Q/KpumS6wY5Q4hUyAWxXx
J1K1jTei+VGUh/0DDx7bLrXFHwnuZmgtunrEhf9NXVuNpcQRtfg1yU4ASocINnEG/mZkbuioT1fK
bioxbG+nFYNvPEmhVEHkaYZKUhy06aQ0OScdKmX0Uc8mrFCxJZLaJ92QUDoTNiYUzVjPQnWE9xlN
5rIIodYOJPkbSIralB9wxDJCMN59LWomffzpREsVMb8qMR60ActA6ymh1wefdCiL5f7aETSxSijB
kEsf7k+GD+n//1Url5XEk4XnEMcvkmIZ9gORCeNcbhaJcy+f5rY7//oYjz2NaVjrY5bpsyJe7fM1
C7UhzVMihww7sldFYoaB6o7eLuH1zbDewo+1/0w86xpC0p5KBuqWQnHzeXdTT9ATg9TiRnw4OVia
VA5FLNXyTLm0AR2YAdX1uRrLAtA1oZbBTtIVGk0d4anEcppPIduYkiGG/7P4UwPUB/DTQRMwkPUI
ikiO1XG5qBBJwHr1nQ4GwHhT6by78eF7kYCqQFs0maUQCpTK0kQJoaeLg1SUdM+RZt6k1aewQcuT
FlpMu1tL5jEYf7C/p3J5VN3LEMWzxJ/nfAEzf7VVW+w2DOjT5PE1YGi2eezE3LX04G5X0uWKCi9V
2AUc45FdjEXHYhFyhl4XgE58QPnV4Bk0S7j/6OQrdZBbhAjaU0Pm+lUDy3a2dLeyZ+Gc0eT7r3sA
U2IvIjlSgpw+p3HC4vATPQa8sHAfc3eB1bFApMcQg6EHOBgn0Qi/1TkVHz50hPe/QXdaDKYF6Q9S
xW9UFsTkAkAQAVt4tHMWK+XGyLjAFDI2Brlw/jKMe1b+DUr7636KL3EJIWR+0eYk+P+h+Q8+Tx9c
blnK8QcjRgd9o7wNWfG59vYwiqmLBHmc550cG+GRsq3mRzKkD8wZYdmVA5FLYmLjJ2OJciFV9Uez
6IZWYEoE8vo0BqsCRfIuc+LJRa/6a+1ekq1JsPmNAgpw6aiATKJqwdAKUFIcacb2TV7mUo1VRIhA
Hv5ETZM6B81XK49B7vB39Zyx/p84T1kwTQ7fhzGh6ushKU36cBLKG5Q5gBXcmvF+Kc01pSxbaFgO
8tIhpWzqmxSSnjpNCG5T+RU2tVuPWAFosQpNs/MtXf8EjVzByZSmSpzmsBxZQWXc0NK0zw3amrGo
iOh7zA/kgF04v+q8bdkRZ3jZ3WLEG17PNrsdSuCj/iXLyIfg0pIzHSN8R8wLU18k8G0zQr1+nz9Y
6MrE8URKcA/RaHoDGy5bO2IzvrnGt6u7dwsOgTZzNNKdaBiWuHB7zBJIWLe5dasyDh2xofeyxGnQ
L7q+nahR577NiodhkNcGC/Is767PH8uYGZdOO2lxk2IUjCvvvux8U6DTSFSiZGbdVKXisTf9c/Bm
0zttzEJamLy7hLFzOLN0emHO4qfUDIeHA4ck6jDSWi9q9UtD5wbMceSsGiuGdk8vHoTVRVc5yJn/
JfTYAzuGeUoP0bols5y4LnMFyzeb/r2AIyJhbnROzKVsn6dodTQBXSSUTISWPHcN94BA9aINpO2u
OdNbA0KZIPFeF7tBqLmIrNfjFCMUF2sOLtctBtdta/rVkeYfzkps6EPmort7wIKNP4nKVrxj3IEJ
0hvje1qI34q49fySvGfOQWoQEhtmUgugZc1JOOTRSMdqyk2fggjxv+jgY5hzH7droPBsPUqsCV1p
Fre3uI+KXpIRskkMffpdB1Jnh6vbhtiNJbj1z8KhP/KS9VFeddKTfm+oowDrz3+0INSOxPMhXAYp
K4LTtGXtInQfecfBRBWAMeYc0E2cA87vrhvC0CWoK4HfLB4zmdFLEFMUSF/IvweKe/uh885Ywc+P
MNn19EvnCnXAz/XFYAtJAg2q6hU+8gsJDTWM77bFNEYRZcJ5zVn8YenOGTmszyTXjOKPwQNCkZXE
HI9UygNngkDOJS47hCZ2zYGR3a+V/ZMN5ktQthL/v1OIZzL08fBJyZnkH3Kcm+KOtquvP0EXFkNi
iSzmoB1OO2DlgYJ1XLm4ffLqBdmNrCWmL89YQorHxc3XZmdLCRyezKBlf4wWCdEF8wnGsfYQPY9K
5cy0+AMZ/1uF6zpe1kWuzulv11qAFDfVpIakbbSDpO0UBm8HwgA8dbUUpqKd0fxhGVnfbnAYg8vb
y/OaKy/uCN3VCoRVpqg+ipY8lP2m4PqKZNeRn0sT26MxlpNttY0k7U/py951aG92NJSPGAdRlJqN
q8z3qmaZWXAMRuWNxEFuaZBfbXZowb+ZlRdKV/wD0etgEcJnvzPS3L/2p/n3PqtrEQtS+3zv9A8I
l4obwnx2dgpB2hs/Lq6cdp4hP+1fJ5CuYW4HlwWWFnU9GGtCoEyUPYiBEAHzlPucjNL+ebhTE7Mf
NdRVSbDjbLhwmqn/afaTNTIsUaehQExYHBYrerLb3N47K3+HDOhgTlUKKDyOywi/qYYdJchMocSG
m+//HFF5Fh4gFBeltkNUpOlMNgG6qquwTkJhNfcCQNTy6OA3txoy8GjI5EL+aL+Yn/F1SVpszGO6
uTXiBP1nj/FsIcryqnPSZXw1XTlUOGz4X5BilmUNgo3v631ALZX/373LzJBZRqB7YftQ3fCKfRVo
e3xlvSzmi0WC3FvS6ozSy3jnDViweMGYBGbugEYWZCNAFG05C5c4wZimAoWXsvI09Pia2WNsaN6O
TCmyWcorMwV2e3qYeGSjCTa4LBT0orYlzAxuvsBl1fXoZbtsVsgwqrr3L1lL6jKRkAZZBoZ1W1hR
tPaS7MULtScIgjkGZd6gNNg3KdAewNT5itgV/NKSakQLc8DtgnhyouX5kNxqWMLu2OdIKf5P3wBy
ar6AxzYBYXpynLAi5LnQF9wWBUaAyXVu0gv2q8gTsR+xd9MC9A0/vs+w9O4LK9NwUXw8vsxccSpo
HThE9tf1b3iuPY7+QcNJP/YB7JmOj7TXjSiV58Sv0LUBwpWLCYavylorv06+BaSxbOmdE9krShgt
V00vkLhHLzrRgkLyaA9o28pejMFcmDvtxVoVVT9uyIme/i1RDUm8ZCbvyWJdL/DKKiff/wHJdewB
vzu0DYXKS8pfOnBQi/wK31QB4eb856dm/kwhK8sJmVLl/Zfalo6RCmTMM0LHpP6KrAaN5+jtI6pw
8UvwYt6etFO5ImYgYSpn2eXfq9q1iA/+Kq3IkXMPxsgcInlmKAYlhRtgFGCL3pWpwl4hZNNYhku4
DTwBs75Ul9ES6Xw5jpnIuS1Or1OtF0oSUPYsw2jtjJRXI/fmwW6itYr/mZJ3K7svOm7k+mlcYgll
kkB0EeV/WGbF0Pqr/rV9bIQUYD5ejy9V/ey8JPYA9onsYKvXi+oafROpZImExEfLGYMUWxWmSbkS
vXme3nTdCsuQLPmfZs/qVJjdCXNLqFLXYuTAcX2DhxKM+xsG/TXbsxy8GFrLW2QwRWRrnc7hKYAe
5mUwDV7cj8Ie/S3T2ajtcUEIpiBa0sMWP0WPUScj/TBhnBXcwvsLv5LFIZYi79cWvTTDbwW77bI6
+4xw1tp1G8hTEMw8ZDDmiV4Bf+ua6IovJS14chXqve2Rm1gjWhkaSKLMT3QP1fvuZXzNSm/zqGcX
T6Bh9wPIRPJO16ORrwZwEC9fJaalDbZql6L7VSy6VQzUDfVGkcHTkhWfDvSEC5dHq50QHGJ3FPHw
z+kb6NEw6HgYxyfRk1GncYN8VsWagZ+i18UJlNpnNtNC0gyvljWFgptsR4Y1XJOqON3e5UjDYQTg
y/Em1uGAe7k7LjVICQJqFD4tIf0HGrLn+ijv6/BOdlkPMNtAdIdyVAe/pEypEZDYV0fg8K+eEZWK
QLiC5/Y7IcNFTRib8SffzIJq4H5fiIqOAjQ49DUbd6jOOgNEKDDXR+1AJHwXoSJ2hIzNDCtWduNv
QCHdTR2sU6ZMkeRCi23k+/hohS9CWLse0qfp7re8jeFzboOsnJXbeVNmaMEDolEQ53kDEk2qQO7j
je7yTVkEUC0Ei3MJEjnbwCj0LQhbBFjTPLpgCzIPoQgc+/ScS83954vthBU67EZJUExVrLwyeZGI
9d1E6eX0ARILPb+VfCn8TyR1e82bFoTohkRlkyaUOs5yRmh1Q/tRAV9trHkQgwWuH6KaG/JjsEwL
1uBiWUWUEthkgHnGCCK9zA8RQsEgi0MvadauxedxlFUPT1DMY3kLtxbVh8dxFRLh+OWqPD7BhvLv
dxaqyTjfSmYaanrFOhwIjvyh1jY0cZ4PgPaBlbP3vXKc0/p4k5hdDvJHbFu93VNL1zrFDTk6uX/3
2ns1uk/3H1UhaI4JdZKIlsqyQ9Ckl4VhMPyztqHnAlhNdBd17KWXesu7KzzaSYa/tz43s8XPoo/M
KU364+7WeMitJl2Fc8vb0uAcJ5ee1S6Gu8hJHdQc7nSXD+q90QSgcfXQC9+xTYoRJ6hSqnbThvBH
mo7haM7LdhEjjDdCg1TYct0+1UJG3WT+4THOuCp3cbzK0StVmyAs9na386bblTkg3MtmPDqTcb/o
4dLw2cfGKHoywqunwuSqcSVO51RNTsNtDMbZDuQPoIuJQPl09ufTkWb2CxXUmOmsJt0+pjvUm0g8
WHkHKPEMk6yZsiD/cuntq62rQH/2luRcbjehqoBgBeSPFqzc6k53Y0X5o98uYQxsNHCyGYu11+Xp
DdPPNyNL2Ix/Ix75ogKcNKADl4vWZVzOGcHKcCmk4EdqunYvjMOyHHocEO2d2iXpctWt2NuiiHr3
imaBBu3P0O4wcfYBplpHYdZzvbeAadxJvKc5R1ZqnzvzVa1aLS/0xnJkJEUhDKJx7QKVV0ITMVgo
EsUvDhq45OTDGkpO/E2fX8S3uOrd8BSty0ljhZxVrl1TSd0sAVsWNCRfw62ES5vMCVEL1eIEHzDj
sflTZaUYSVBDVoAwDnHr7NLBUF0ux/1fTr6XUMBkXCzTCtI4/eh4u+eWBauFXUzSO3muWtKi6COF
D0OUzQ2uR+LOb+vVKGKyYcOwDEK58V2LrVZqJ0zvHHSEN1vmzA9q5ssDRmGRBBt10VKd9+e8fudJ
a5ZC1+fCOiLyU/cq2OAAjT05WY/T/nIeR+7Yy4ZNOXBifNKmuAbUIubsCp1obEBHkF/k26l8ZoH3
jO0F0xaxzpQEn3l9mDFEArSCbtflBY6jUyesy/i0z3EkVyWA8DpkD6HQdIVsM2+krh0YMzSEG9EX
N4lVRkqeGi8OKFQV2VNHFEnCZ/MLdM+b+LMb0XwGJmjtDvwA69N6WW5zO7dt/F7pxNJcdUvL79Sh
YO8bYGyBiCU9CU1xYV7L6ygwZUdkEM+QjqvG+dcwziXsvHeQ8HGMeJydw5ldAzCr7mYvvHKxK0mb
8MHKSB1/mEs1N3gO+WV6vs1Sn2gEanpVywUoIE574VusQhJeIwP0XDU+nJq/UG0X0mWgjqHJ40va
3jtoZs/LL2mWKpXRc5tHOaPBw2QiN0LO+8p0ACIezW3VIjNQy42Hi6yG3VuyRmMm8d8NruPUPD1i
ASo6osIs3rtkVXlCsqhTkjMGD6moAi+7uTltqesBR2vrsLPZBPgBmAD51dceuivq+F+6IAmeNzHK
DYVdBRYcu+qGK0Pox/n3K/oDVb41jGr9whKCMi+1Z7W2JdtIzXfA+rk+iF6XNVqNH2dmS8DdoDAH
CvYxt1xxQ11Nsb+MG8o7K7bxfgGkShp9U5huBpiNDAy4SoiO6ph3bTDsDRnSHbE7ocwvSdjluI6C
2uHOTja4Ge31tgIIzxCDaJA18MI/9L4/X4etZhqO9j92oEPOg4/7agOehnfYKu5sLeQO61YTFJ7g
+i90Fn0Jl5DpJFXdLibqzdaQlDtzc83/G+2A8ArQRU20BSYZkvx0SmmpRP3gTXbpgXyHHs+7MrK6
LKfG1sm8ny4ydqTC5MCQBMgcNC3uRknW0rKcTbQfwt0DG6424z9JCQxg1BPVZQoa3TsdeDY1oig6
Xc61M83Eo4KzRdGPiYtTEhBmbhO2wm584CQCeurzOJ9u5ZF2hwA0Mv8F4J71izxRvT+6M0DFuxCS
zoLGmeLl38LdRG9rkcClvnB5lUCCLn+32VoLwugoAg91i1oH5cXWLIWbGNDFke5o27VON+nfsFb0
3kQ+rqit4EzPfF7QBpXJ33KIUENwuWGOaHT+PSEyamyQ3DAi6/Pcz7YHMxox2ko5y3fwi+57PbHy
PYu0KLEI/gZNH2haPsYzTuWnw1u4DBhDYK4OsLSqvq0/SslsaQvXttrCGuhcfiqyXqH4Qh6gCO3e
Iv4yWuU/mAvrtMCUP1iNGE4IRKvJiR6YopUeDZy0wVAXeSDOQpzHEHKu9QEdS/NUiA3xM5cVB7fX
VWNUMIkQ8Q1agGZzCKHPV8aChGJOtw2htzy/HXpx3E4bZjG1a6TKTQ8ho/cqf+trgg11C7IeA1kh
mnXualAYMrQmBz+2vo8nCv+h2qStfdvZMBQGoGjIzR9wNtCJfkMiKYP+DiCc3HIntjiyzpJzPu1j
qjZgi2jsTn/hMdHoA90PBZeoERoeyjrvRueBopNkkeY7VQHiAqvUYBmCXxhL9PXTr/30P8DwdpEV
LJKgNPuHbi5riUxcliHO9HUKj55UNOlYmRmCMpBnfQvq3GokYjzEm4W3/qLgtnSUFMOj+/mD0Mwg
wsAK0m5iDaxpeL0fX4MobnkQD5FM5pXU1vz2nAb49W2Pw1eYsK1zWT4BCyYAFON0FbQyqQN4FSlJ
xRBZL3XpsxU59OYIN8YKWdbSvuJuSLyk+M20JtsR53pkg5GIqglPV4a1Y0X6Ky+8Dlqf9Oxqkbdg
CCCDlqPmZNxPaELJouCORdMO7Xtmo7+6XZOVWZ1g8P+rpzzigWltxMSC8CjV4QuOnmHG1K+IrxhM
yDk36olKI9h1s5HncFy62FYGfFda/a6q/thIRgsa1MZt5SFNHv6OImTtA925msvvrvypPq9i3gd1
Dyl8xRRVNStqwzzdOBEdCsqb7PPggUUQYkdOc3WONVW34gjs9Ez0AWVp1MIMJzThk48TPc0ZgnAA
rYYm2vW8wBtifeezZC1ymUkEEzUNg9BQ+e4/Tp2mKFLpszKdmt/RzAkBO1uAXfxdl5y6F7HSr7TF
WZOZ7PsgS6tBfoZx/ImRafmwN7mtdPMIt61gZbOEHq01QdSyh67lh8D+IN5VQqxEk/5hd1McV5bl
3pb+yAxRVtzs82a8iPwgy5SGSE0mH1EtEafOJpnkg+rwThU+Vtyu4z1C+EiYC0JGg63HJZbn6ED1
OEPNEtEsfN9Gj1ppLC+xsYoN/S+6knJ0qRZnsC6114deyIMprWjREy2XJDxxsuragUQQAgcy3fbW
DOl8l4zo4HYqFi5GkdAd1KgmDR+WIQpp2Fsz7eN5BuvXX467xUSDqplxyIvHpziDGG+KcifZzC6X
yoBqswksE0R1/101WKvVoeoC/zkr3sIJmPTUZlwPpMtlZlGqIMqZmF8H2jr0X56v1ZMIbjdBBzy7
Z1dZdbqA9GYOlqybKR6Ya9iUXZ2UMSYw18YEGi5vqnXAA/fTMKhXdanILpFbeVpI2RDDvxAYrxcT
A8WQ8NXNN/D0mwfDvu+i3I4VB+pCPvOw5EoCcIUZLGSCJcYdndJs9WqENNrczg677VZsS/ylDsxL
j0c1F9OMflGu1nUcxuSknKDDNGt6laKpKJmi4hOQxodzQGAwghQ8f6FQUasRTyqoFvjwWCUnvGFi
W37kqUSDOxIYbZx7E+nYSaXJfBD/67xnxAin9SHhNHReUL+R0te/d8DTSBK5SrfiWxwnG4wVjA8a
jIpqlfI9/xdNBpl37qt4RwEkKqxC+6UzPWGudKUCitirLdy2jdPqN23sfgJ7SznuNSGgEkG86rAR
QsuGQ7YLMLCrR/gnFwmUWBejZM+9mzJY9P/xmMYdCGNDwwHoydKKWZILv8aEebtjMHIaLJe7mZmw
AztfAX7JXwkquYFz62yhb7fCebkmvOzqDk9LUkUPcu1Twl2MWij2tkMKZYVdOdMFImwNG+qYPAC4
sKxuByqlAiUH38zzzcYfrxDPqS4iiuHWJrj6ilZCHzfOs5gCm8I3PgIfu+MEkgaT4bRumwdNJwLy
nFW2Q8CTHycrTGspbHvPqZegSG98w3TqIJDIkxK7vCtWnyMRInOwhSHj/xZqQ70ALGmhK+lDgsOH
MZeGlfiHGqUQF7lPtC8eacYih2gG+d2VtkJPo+H062bJ2cgbAh0AjPBANuProzmzgOwHrVT/a12Y
LgsWN8jfaLn0ANVscZ5KA9eKUDnVfqK3a6hbBBiEij0Z3PQQxwTDDfdIMBf7XtDvnMqH6Pk3e0oN
6puYjbfLOdPTDXZBaKyNphwqgcZDN08crqN2ktVA2Icuqxr3UAHyR8QVjsnBHM8+pRXb+hBX44AB
MP5ZYQ36hv501XLqyMvPaOsDTDF452SQ+A7VdSilPeArEAQncxAAAkeh48bosvNYOLiQYQCFFRCV
KnnQuHgNXfoS8030YBugvsJb/p9YHVrNSFpE3LAWvlX7RL0Vps/TATKO49K3tEY8Nw9G7rgMhUvD
5W0mO2Yxc5PvGIR41rWfYKpetjjjVCLxYBodkc95sqgvJd+VdGTbvjlLj3rAHieI9LdGN7ChrmA0
U5pm5THJAY7INKXPtKIKeyp9JRv4xYHrU4OZcVx7zVlTswWMkvUzwHQEnKzcu8lbnenHwQJEwhBs
SCGZXTIASDDoEM61LXjvxyK7PlpG4TcNoBNsSlVxtkjH/UZpWjqPnzg99Ga9NT+H1NvNLbU4roIT
h0WVHpCvby/m7tIe7oHphA7x9bgVd42rkSVC1TPqDTjo3t3YLz2lvp8jCjiUROcOBnu6oKzzBPLK
cggAtZZPXrx0pkdgm3Sxg+XqHOXZEoM6T5hzb6XeJo4cjz30JxkWqZUJi0JF4IAuU3uRCjUO7bOP
hABI123ksKOP1qbEEY+1gYvenns8mNPwZCQUPinAjbMNJ1x8DRtJFo7V++HL6fIkkOltvjiV6Nlg
7fs8rp2Ylze56jU0GGodxvd8HQMfhloY31jA3+GMvhSM7ZKitwuSX96caP5ykyOf7cZtrUnIue3j
WSWS5gEt8Ge5ZqqlJwBMKG4VQmpBhZNq65M/nIQRDtwMeeLuYESznnFPiEVH3jo5rS9/IMid27+Z
n6N08bO9SGMUXJ2f3g3Unv4iTWNmJD68wqhJczhT0PU1am2k1Q9bl/vj6qbQOuNCzFj1vNg7hd6i
Tmv81shLox3gfCT2hC/bMNR7fT88j1zSStk41Sbca3/xA9YTVNxeQOhSyLYv3mGN5cw9oB1CcWhu
SJbSs+JRnK8vLV2/m0WyctIa6RUwwwmDvqCALtzdOsza3AY/da3LULBKyPCV6017hmxOj5RxaMCj
Q4Neb83gtvutnToVOjtMr4rpU8YapK7EKXW1WvjuJZB2nBgn3XMTd8ZYtklT0bMpYjmIcqEA4Vn+
saY6aSWVB8FQG6A3KY5ZxsGLFUw/DwE9c7fplXM5e0kBcxjrScX3Jjg0N/3A9T1o/uns/6udokNW
vanIhSoEWNqIjTsLkWUneb/7i487mPDoKfQ+/DjADgGzMryYwGbQKpWtgFucByNUTLZyNclQYQ+0
jgJorQfVO4nNoluEUNmCD1ZmLnwdN2j+Gizv8WZdlGUAQL41B/onZWNpCfD+5SqaxkNa+2ZyNM2E
I2JZBrv77YtO57O0vl3/sbTg19JMG28/D58OMwWw/6bjlT59y08X2b1x+fOFVdzQjjacK2lKgbYL
bM69LoyIK0gSetFIQnb64TBlp65/mzMCgRnPchivKhj1qtktmGX5oWA6AX/mRDlQxyN/XJBWFbH/
lt9dAlW4chHYw2GNjz2is3QNPntm3IGwnuHLRiNbOccyqhQ1lz3OoJcpPk/ifFhSZ7zqyGkSvoJ2
7+arBWo2THEfLlz4Ppai+Xi5i1GAfK3Gnha+1gGSgntTEyh6gG1Tm2p6EXXhPOqLbVB0Z1iSQ02h
UKQqMTtCqt3oWHvSqniYd53TrYG6O+FXrtCR40SYuAIsxtAS2YK8LYXk351jW865JuuK/jwhed4c
AtZGbaDPbL5o9ZbdIJptEuEd9CAT1C3AuYdrgeJyZ3pvHNdqCN4QTVDuDbXLHU9WX5eUYk3V125D
jCL2D+Ysnqv2yxHIJAZfTT33fdWuKzb7tf8GGwCdefbbbXp7CqNOZUf3OA4+Q4xdDtxWrtBMzvxp
3VZSVSAwHFmxO5/e6aCSYLI52ltc8+4L8FuHJjO7P6KATlE0EyPAzJ8dLfoMMdrcdx8Hn8OH+acz
V5UhWKqkfgSJsaWoeKrIxoFDCqTY1NuTq3/I/6ezg2fxx2N7bhB+e3erKEzGoycrR0DaxqTVrLIj
A4NvCvjwW9RpUGiz0iRScBrIrhrijHdvHl2D1juwi8nDLw7kgsx1WV11llMKesNilRiRgVpQaGdB
vBAX2EzPeQLoZY8yxjph9hDyMWjaj7LDCyg0OnTnQN9LH+LGUYWQGwFrcRTUg970GXg4/kdU2sRr
XFSGXORYRjyUZBMlYSBBD34+Pzv+UkAOSesJz0ikaDrC0+bZoYDfQP44fL4VtxJnm6z0OM4Uqxtx
7Y8NRZKTNV5m228k8mnGxEOfqNfMSb1HI9XeWCVLcipe1C/I/vYMczSKnwB6/ajzIznxi2519WXR
yP8hptkGHPPw0HsivMKDfDn4Z0iW8gCl41/Y8OOxEkFS8Y/5I5QltdFN0Fg07+0uS+DkpPS4C+D0
vDcHU2NVCtPEwQFicGj4B1BnDfq3ahp70hhEWuk5G3MldXjlkwI77ujEEtkjP3ZetWjRnWfHbBOb
FtiCYa7SBS2GYnhtAB3B+9dXGiRbQ0dZInVkxu52ZMfRwUtjWSgbXrS4vpgoFzBQR81TvZGcOET3
8aOvQzi+lLvlMS2TuXTXe+AgpHxMjpl2iuSQ8MtaWfUIdnBRDAhr83DS6pg+uRBbqv4KGvG4iweC
S4LaLfk/tqvQ7aQF1kfFeqgU/yJHGo6X3JFW3EnwSvn0BgkzoWO856tjOUzhNmHM5oyMxxmllRvF
OVfYV9lJHeEWGpFW+wCHuKFJohw4GPp5JjhNoCjqnAu6RcK2AXZcVua9BSxFx0f9e/ERPkdmckHG
ZQPljMTqp6NyvThl7c1su6K4q02Ci2QCcdreJlieXoZGni1ucbT+1ZGPUs9SfrthqlVsc/dR4bnG
bXT//zSol0hahPWfe5F8DWxMsJ00hxn1OIaBosTOzkgxShe9v2MSd7U1MNRqaJqVro/w8vFZiZJH
1owbpk1qoqspnyDv4WBG9+/rDgo30fAklbBi4A8zExw04rZ8OsuP7fuTFrc4QTVZe+II1SGNL1uV
uYbRR/n3HFsRVv6fXpWMIGJRFgNXBZkyi7wp91KbTYwMPjJX7kxNL5CPdg8o/ANJ0OpukNncAxbR
5Qn7frffcmVLMYcNtdA9gqYXNseTBQthugK5KRfU0UT9y7Pe7GXyaqMRqtJsAwLLNbQ7UlSq+sy7
hcWxeNjNP5/lTUlKNf49ZYC1SoUSkJNjg3p4T9DrTQOqEdLNbVY/M9e7HG++isTDhcb1ObK4XxG8
Mr8aJXaQs2ubhMfflwWVbXP3Gxy4S89EXJKR2Ct7Dq+f4rnSk0KGox0OS/RFDhDUPoQbtXloozZ3
6x+qk+kD8jBl9wIj2yCu/ligXbfC8jKQb5PtyN4JH4MVqrwooyWZYaZtH2Bb3RMdgfZkgXGbC5mc
IeNaoXsaqfBkt3g9tlPU8SqwS/6lsmHKZIFl4u1J8Th9Jg+JT+dC0qUKpperhwq8B5opVdN4r0SC
qFm7AIy81OTRPDIFIpaPHCoUVPqjl0P7Yn3HhUxn+3EhTACfwERLgZkSUcXnW7NlB0kpDVXkVulL
q7hqDVL7CArTp0Dn61syK8OjyCu/ID0/d4oYsz02k8lg692Ps10PcL6MKQityTDP5iMotjJAhIIr
s//mE/mV08u7cZJBhKmPO4Xhdw1q1qBgu+Xx8lQz8LQ3uCNVmTXbU5BVBGEXoPouZbnhF44GN/DW
OmAttUhWgKaebNsFspEjLERhveR2h4GYJQramaGcES9u7zNzVZeYYfL1qJFP1FmRlQp+X46E4qqK
vA0V4nVYX7YGzPZVA5mGl091pkiCk6Cw43lSUe2BPBwlHreDxz8i431Wxsv3hDwkt/naP+b9MzJK
YqFIqHfY5nVKEdZ5zJ1fGqFmJh5GtMbdSLIyxoCaPorns7x+uXAruZamAybvthcBuh/mQPlNpyjS
aNH/jMnAziK5UEPkIWTTvsyXj/WA8mLMDEL42ZwG813Ye8PtdehnzGkFwOiHMmVCjcKRXNwzbTaJ
pDaZZCYGe6SFv1lLj9vb76UYCn/Hwoo+PpcclfEQJt2YW3qP5bQcvN4fCUO2ivV3w2QvqqII6NZL
RcPzOF/S6FugELUBLa2Y0Kz3O5pfLnaPLRYt7AqgIsLuOscpTJMm5eUkrz8gnLK5L/z9CnSYfeVq
GQtAPtrvFKAbVjkIsOXwBOvw/wbfIbBUcbZShkiv0OyGS5UwIhP6hiAh04HaxAFtf51gWj8HMAOV
22+0wt8krbfhRsoMlTQ6cDLPiUOx53F3WVslRK25pe2qYaC8ZkjTiuavqhisqCc7YvnDw3vjOpm5
aMNqs3XG7sTjBNPNKqoIR4sf8HQjALZecUVL9ZdY7pdcKdDjjo18N7egpZNLpOfjnydfH0qWvtuN
tPDLa/U77PPtoxQn5E2uYysiArGLVYNewA3wn9J26SOFqDnGqIryZbuh8j2BXqMnCK3m9aq8Aa+K
F4uR1IMYgXhH26tKxK4DUHqck0jXc+tRn1HxkwwTyr/F0KutW70ljZ/BmF8/HL14NxSVSfE4WZlm
vpX49tzfc4WZQT2Bb2vT3Qx0+eZM34hzxqZrPPT2JWnUptrxM0Z7y93ISJidKJO0O2jHUCO/6uiL
RxrfAOEDqkkqbtNj1urVRr6/ZmzUzCXQsCum4apfWfl1ZJgGBmyiIIx8tOZCuldw5To5buDkaaY7
a1VV04L2whr5vVZDv2PlXgpIFPjgpVn2RWLAnXqUJNVEj8xCNhI7/ma6JAfz4+elYTzNScAjvgwo
9+iCEd2Bw+MSfbOiPGLOlic+LLVIpDcqunHk3F1/9QUKEXngdgKEg776VYDxWcPfs5qDbHy+XrH0
rwif8K7RdCM/t6tK0qo1me4ZL+ViFYcc4DxHYZGiVwEQMNRACwpI6jYzKIL7LVkbtAUq9Pgvm4Jy
CwnWQ5NWLykDJyWckksOWRzGlaSFLfoiGuAj51tGw8vzqLHvu9WvY7HTwV7fMjVPX1ssYbk2gd4o
9TteM56ytKmPE/j1wCScxeaNfeJC3bQkZcypMiPsryYALk/WizzCqg3z7+6R73h/DhWreOvmOGc3
YA2EOM1AKzCy/1Df0Qcks0KHeEqaV8SPwtiNaMX+Ll5vsQSThMQIehhqggwRbTNClBAudlAAuXHP
P8AicrZuR7EY8b8wZTIIrGp6hPuXLE0VUpUnbLqDYOqvrfzkTH7JQsr2H1pmBIMfQ0qk1CyVYgGJ
izicLIPOCFUvyMiZvgddFCjkgBp5tla6/A0TbMLwATYSDtpYCr1Bgn0xY0d3mYg6THqmIp5A7faI
iOLiuMrhK/KxbE4mblqeaXtR3JC8v5IYSOKdk2uZnf2p+bH9c9mtp4XYEsUwRWbzUg50mRMOB9Y2
LEV7zV35jV3BYZ5saws8+5hT2EMRTYSKYLNHsUCIdf/yhRyPXsm0B0Hk8pW6YKi7kw/0voE4ZNbH
MAC+phpELU6IpHWNiBlskpeSohUObGjJyPj28va8ki4HEpBXI8LlRXBAFbqXdOhBeuqoStIiyvA7
Vu5B7woT6Uq6PY1WhE5cpY/iGMX8unvVrin+S87wYGxfCLWkx+Z6VbEsgsp7tUDsmQmMOYepOyyT
MOA48+WnI/cjLlQdQGei2ECWibcgyTTkl87QT5rjh106RhAKGkydHJV6jvY4B1vrcs8sWTz8DXRT
1n6PIQ2BNP2XRqMZ8tJV3LkPkrdKsjW8epQUyOPza+Oi9+RKERq+4qvIuj/3oCnwL8FV7w3f6Maq
z2mnSPg1FnUNHeVyLNvnd6am9rYZs+E6vL26iGAA4bk7Wh9IqvRG6Bfo1OcVviPDi+XcBoyt4rlV
NfxG0St8Jqs1U90ysENichjl5NHo8y6pRPV0Grz6JNXwz7zThD1FRd2bsEEHw3Rjx4Gu+GbnRLZA
AVVqT4MbyHEzJdv7h8uxgc3gWS0Hic7txe0+7rKVtZvy+EEOHkpZxUNUKXzUNCSFUsTqcAh6Kb7p
O94d9CqOciOKLN2PuSOGeO0/mM3W97rthfhR1vIeLifcEPRllirZe3PdtyNTycTgo/bqxPsqggeU
oWg+nNCMFJMYFct/CuOyqnQNJ5P4tHnB07y4YInrTePY7qP5Zbq595VZ7tFzvrR9DsmjKkEKtFKx
IU8BeO5Nie7O8iF2FJ09F/CQn3sqJBp3Qp+M5wR/a2WUCwUJfxAQ+WAAKc7mggPSBBdVskeWIR+q
2Sm5lb9DVM71eRGCkNufS/pcOc5iSSIgQK8kF+m/BRKxBqMgp3DwD+OtD6QmQ5QiJAhT7BduwvH1
bLePmZmkRMTg6kYcLBDsbm3m/UFfcj0tTchkH5D8/w1VRyC0VK3Dlh6YZdXMQ3PWF5kzDojQUCIF
VWaKrpkxcgA6y8zBndzujOgIF/sHQu9x+xU/pE3+fpAnmEyazfDbn37MZwW2rjufoMYuG2A+iQfY
96rnkFWUaHzvn/UOvsdZjlLBBPqS2zPpgarqqkjtWUrv1SObXtiNRObEHUBSdb08FKwO1qJ0x2/5
ikbf4x8ejPeOqRKd/bEQNjCQ7i0NOjpXUZwxi5uzIPnd/E9w9Ob8AsESiY3WE7GVxf+kIj0Zlos+
z4WMVxMzxsrbIFn4uxszO/rvMoNK/Fv2LK1zJs55xidahDAyUqh38Fv5JYuQjj5XZLXSFJ+2TUU8
gh4UDsd7X21EFltWNvz/pz6rQDunQndza2rqZFZl9bQKH0EdtyrKm2lY44kg/nGjfJXotCdkzvI1
GZrLqsi/UqcsRDO1PgsOz6V0tCTJixJvNuuT8KQeQxUaWLxv2cHD4yH7I/857zW2cK3yV/lpQp6v
6cHFCGt+WnboPtqOPmbv1UlZUw97NNEolBluAY59TY9JCKi/9ynNK3lTcv/csMdF9PYviMObTmgL
Q1Hvxqrog86aGX08NRPP3QsDAJphfKmcL1eQgIfxgU3xQa/oeSnrj8vzQOFUwck4QCyX1vCyqDUM
COyxB0vLTCxzSQrc2Uaz4INEA2fbVtN+3gaGJ0YuNOBZsHCUDVy+cNOQN3wI92rsZ5WuTXBBPNWR
FGRYoFKAc3JNw9HRM0n9yTRapEvUHnWNuE2Iy8Ro7RfSuGxo6wiIKrVwnc15wDEZ0CtuZv/kyQaX
r/daOYOYaNFDgQ4U0o2xsNpbkLA8QIs1bX6lE4rMaELi/oCaUaZVHekdgYyQfDswnvduItEq0SCQ
6XNEst+V+u+GrbONc3Kwh1wW/zwwLvvgL7H+Z8lSz4JSVpHke7dL0NGtASa2zxSyR3Toa99Kado+
S65pCjlqyMYZco8Sa2OSWtyYGXH5TyUx5jzCCLkUaipKLg3p9T/26uVPKmmmpg5XSG/e0yKKVxr5
4kvp6rnpAWiLF/oDL3+jA9ZzhO1BlXpDyK9bd1HN8he4Gim0hBWY/NwvSJnvUzFJuhQGM5uNhECR
FAYsVBerMsM0schFuQ7fcLt3IQRKlp9vTtex8jFPp8m3U4Hj6PonoE46p2NqSR4seYxQAPbYDmCF
Eb/VQzH/l79fWYZikTYkqLHKht04CFIr/zNhh2YwsW3oCpnGxAYgZv+NSVZZe9tU2agPaf+BDR7w
reqgm/72xKGoZlN1ykSG1uOAKrate0xDnDhpSgFxNI70a5SuMN4tihasG6Yq20wx15I/iKaj5MUP
UTkI8QNFxr3TD6td8/gW2VKgUIAEIf+uzed1drnqzpqmusLP4aF0DYcU/Dn++ExmZMFQtiFAL/C1
5m/2jKOeU56QDCZXWQpH1xRt+wxEVoBP7V+OQSiX5rVBxtTUD0riprIf1KDmWm4CQpvo1Wi9dPri
/F2D6MAk+kuYxbxitlPNhbTiJzRhk9eNXIERFQn/xXV1uGtPMSyl5LRb30q3Gjv3BXjKZzZUFrCg
7NJicp9YlNDMbDJa5xxb2YQdiwBWg4NZaATriFG8mZ9J6Q6OTrsZpROm7kcA7+A+eQ3Zerl3u68D
iSKa5jvvS5Cn2AiSyTSMEqCCHOxshwFby3pSHaB7VErs/uNc5eLy4szzhtz25cmX5al85emISmYN
sFBgS0YmhCzVsiwaszscVsubuEcyqEMzZGapORIlqZF1MD6sc/mPDAujWSRoqggxeiDU6syEYwgD
TqwoaOyGTtY1SqwULm4g+rxKNL4yvExoQKn847QTXFkh5/YAxnKtRBKb78x5fndHBF9AXWMf0XlB
U6GxodtjIhzyWCGAkKNKdTc0y//L9ecSDqoAj+eK+/UfbBuRBAGBjJA3Ux3+QOFFfs/450DrqH8S
ERg7/lqkNFr4hZCf78CEWO9WvCtNsMiFCAmPpFr+6JgCNyG2qkPYPjtTSqj19juRphRD1Mqe57V1
YTv0at63xuOOaA30JyhbOMbWHRqRGdEYd6vEIQtCwPKFDxyMYjTJnP3u6dQB8xf7f1W8HnLf55JT
ZpvT8Q3M3HyO/Iy1iNfhAm6//VntvIQYozU+kjxE4s+XZtd3hIn/MbqwCb99oTQGK7VCgV7eJ89m
TeNA5M6xVdESNgMPQfevklLo28VFOUc+uWHy6//ye3K1JwltiozlwwP5ScyKQKMQjuH7uADUHX/g
UzexzeDkXHUSXdRapwgPtPZBWx8znohAl2Dz+gHXm9Xe3FBgxA56Kl7YM6ErvUwWxC9m9TT2rObs
Bv4MX5Odxw2qOh+6g1Nh+9ME7LqFGYW708j1KPDGvcgnI0d6ftX5SluHAnOZhjq8tbwLxw6DxhSc
uCeQoy8tJTKDqKfIBfR5o9nJk2Hz7RnTvc339xwljes5v0l+4WHABuc3Uxt/5aZytbgm+KxRtKLX
a8UdmAqoNXauhcSHgD6BOzuAfcc77agu4Avq2xtxOxtbpufTYOyKrIMiLgUzeuvQ05UKn1CkRmta
0/fw+NOz3xTmpbwFMuFM1o8O6/r508WEO+pD8x+79KIk4UMsMMR96myEgt9HwGxez70mAuPP5OYQ
1p7oNj2XyKp6cB9WwR7s8rqQeSYggJyrJz//IGFz0fYWcrDNdCzAhNlaQ3N4iiiwmh8g2z1Bv0zZ
yMRsMHtuhAms421gQzk0LVChReDF3rJeh9YXuZrMQxfx+L0l+lSda3/1St0uB3cWtcmr/TDr0Vk2
X5hJNUstLlGoD74L95fOsiLCugt7RpJqFSC2wNyRRoQXn797bC/Jn0hUfCCUIaVNO7BGqtxt2uuh
3qZrPHdXrbLH5/PURu+nMKBqxi/gbn9HiWOtCnaqri1O9AWOu9q0UeSMRGECC8iqQ5njhcOSHnKN
C+tC1rV3gJrJ2pSEBm/PmuzJgYdZdd7EmVOgKSZ3UlmXKDYUhLTP9Qr0j9xXIsZNzg7bShYsLjFl
k5ES+0P4m8CVKN3q2PDCIE1kEB6jGlcUiAipgcetAQP0bm8Gj2lIolwf+9ctHHQr8vaONovFi96h
bjBTxK5MtsB7j+voC9DsQQUm1rouQSmvc8Q31l9UiytBahObUHNE/+NR4DIkaPw6tN8U6iyCeJNt
hB+hU+kEDG2SlsD7jVJrzVZagofVr+oI5uUoEFgRSUG5ydGC9SAI/SyAaQxQJM95etDoG92jHhGs
UqSuuczitsXFgrjzbxHsolq7fdXIZjBNtw5cwhXeFgnJYe83rvpNgo9xMKgiHXJauN/KEKKzSpNP
jPuRW4sA62uIogc6nvppLJLymxB0QgXJAGop6i4fx4h7n5IwUS7SBRL4/iizLBj7x99yIFAW2e9Y
z0S+rU5KR4BfEAFY0owN+YLydzNElybGOgFykneUlMAGJdmqlzXhrgDToL2ZdJQs86efU4zDDaaj
5YWsoJG3nhzTexr24oneBJaIrszfe+ST7/uAVTFbq0jRb2OcdREs05kUBLUH6CFNX6VJchG2m6oD
2zZzX3XGlGCSG0nMQmsODsfZTwy68zphgBhuUiwEJJ9D9xhWQuxWfe+MLYzUTvXHrA1noVCuu3SO
JVRZfM3muttuw8gDhLgrunWODP9Kltl6P4RzDyO1tDGbFCu2kDna3sBelHq4nLkbz1rbfkNCH/OA
EcItZO/FDGVTpO6YCQ249FGdb5qDHXxNXrEFITkvBF+GGWzjQ9sbrqWiUydaHByNuToE/OqYRfU4
Z6gnKOJI7GlANBVOyV4DyFzYjdXBse+FN99SEGW2eeiq8RQzSWiht29/WlNRNLLGUI470bUL45mQ
YZc8YV4eysS7Ng8qLLoO8wp70Jcc7PQitlGW/RjE2HxlKh6gvDxyGwkaiZp7a4eLy3YwrifkPNb7
qia77KVOyXbX6aXRXjZ71qWUdqJ62oCvFzXRnK2MakdARhiiSBRtxNdeHegH8ft5wb5F8IVgPq0V
6Kjv0BTb3k+A2jafU5fSFStYTVrRgSJxXD8ZjJkC0rItqRL+EwOz9zfpMLivKN3BZFKr3hy17Rhk
paybQB6rORSlz54sfP0L805NeJixlJ3oKMEgiwW/7VMDQHkYDLcKPHs9hQkPpIPUwNxfUxOMCd8Y
cpRrZNnK9/iOsjVMdOwzivrie59BLpemcugrQrDm+DvJVAhcNpBl/6WFH7KywCBh6n8/nl5n+cWJ
XADJLLhvz4yLVigJs9emGTj+fSQSsgeWxlN6Or/5ag8qzRKkihaY0iMx91qxP8EhQToTlWxTBmwA
aebp+6ldZ041HeGUVWeDZor+qvqu5TbRy9eSxvGNclI1zrdxvczb3qAsoIfDmZFOCN0tYOyQJUcU
9oa9DpmL/mF66nYqQwH66/y6p6DQiBETtgVAfbq5GGx3e7vJ8gHLLo9MPp0cqM+8u/vttLST5hfG
q0N8+CwdDvZ0fDp9tcyqyaksbkNooUZGdAMUP5sHGSFRvWru0ALiuMc5MoStMIdyNoynSYqlR9/z
4JAN6pQMh2taeAf2o9cmxm550irS5Z2JNqGcjOz9CNY41zCNWpqs+fT0YNIU1wPcLejGWLDoaG3Y
9lPsbnu+sEkqXTGklU29CGW7v7ukiHoBsDSSKkBqGHqdc+qLMHJVxHux6HTDEtYTL1ebuWwgZj9Y
qTY1Z2dx+5ax9Gtk3Odka6BdHAvHBZHbrVAxtQtxtaPaLh1aLaMtFG5t/84EeCFrqcC2ekooYb8q
ABDcsUct1GogqryKLgRz7aDvxt2nfj5uuo7GW8g7FocEPsxveZqiqr+yogWiRLspP6Nmqlmrlaed
1AmzR4R/MB+0zTnO8iN1Tl/2rWcIM1BkaDsW3ON1rwN4SuD+DXuLC4CpPcQUZ3KiAgdsCgsQyDfp
HmeBIQ4qyuumVN0ndSJnoR7tIHMWgeCofaIdFSJr9c4wLGPC8PQa6ocXFjkFVR5Vv7r31OK6e5X+
KF7A4o5tvrQkOFB5lfO8rV8dvPNijAwLymZSjSU2f5ZhCI8nCmd+s8zG3NqPiFdMSDNOq/OHMYMC
SynkACnu/QC3apSq76YWrNr7fyTsCad53sldkyc55U0dArg4GnzFhm/qE4J7GZ7txyRLq5mRtgCK
joT8/eQJcLp9Q3ieyRVFy8iJoSOyex0AlJf4EnjcnMKKWoJ1s07J0k+GLf1d+mPDhdy66Dj2xfHI
f5MC8mlMknaLGCBBc0NxYG2Q5FmruSijderU1qCXZ5grKShK95TAdhIWNJGHUoJH4857823oNkB3
o9nTH6PseZjmO+7ij7exkL7NW88uB6Tkr0x/GhVwnR8iVbmRu3+uGrb08lAp2XaLRpY8MxPZ/+Et
svxWM/H0cKom1Bg6c/QjR/y8HUaXAHeSFV/69MgpLAnRx82+h/oaQP1glsBAu0R0QXLsL9hZwZma
G4Q6COcPvIflJN8mi/TfnC3WT8a3Zqf/ifmBs5jDuvMfYaaoQjBRLnUnOSVZRfYf80tnf5dGdP0U
ZeOOHmtIPU4XF+9MhQ6e4JoN1bZIFSpTOUP5JGH0szevte5n6m59RTj0MwmZa24m2qsvvwn5F9sX
Zn777Ufxf0h2Z1X1weafuJ72tfGSwbONHilQfRR3aN6CC+Nre7RLC4wa8S350YoDm6wZyzmClGlZ
KMaSLolqo/slyBvSpxoWt5TnUp+VIRCn4xA8FMjwWT39ypAkFjnp1MRj2SSy26Bl/OnuMi+pz7mK
g1RFRD6gOBUERVD0tJAsMclISa5W7StT6PeLxVFWZfuaLTVoxfmtXRo3E/cYEmINt2C650Gnb/Ez
oaHMLhonstpHVBgrsgGmTJwy12RN0neZi6ABwCFM8JH7mVsrY5GzHUIn2oOJPUV4Ibef/rS7UqOG
6aPE04Ecms3pY4JhmLCNaychL25vEeICEMmq7C7POywzpn5NYOiGrSvRJYtPVtw2/iE/XQAu1GSs
ZtFXGYAWf+EQlrmO2qP04zuZ83JpbHqWoesaja8OOeqZo/4/9+sraJ5g/HZr40hSdSz4VHXix+Is
GbikXSP5LN3pQ/Bhp0mwuvQlqP/Sd6J6Q+kQG2gtpnkhLbIijlqSfbwP6EYKJwThFtfc8NHbY74y
B2l2F8dqNcLkeh8BV1VB0R5SFg7voN+4AlsS5Qu0eeaJ9T18SpdhhJfMAcBhjQd7YQf54kmZ35na
WBSeaBHYXKIh3QiBmhKgLv1P+1sdu6PnX03V1gd5nvKUjX5L7IIqKRH0xEyai6x2k5Upd40IXh3f
9g9mrpliiS7VyioXvMMw1kM+++eY+U0G/PcZaVeH4803g7f9Jii2aS2SHAbRV92F1tk2PctjbNqp
qWlEyzNzxrWSIUGVuqnz5x7qd3UbIfLwSzNq+whvR7qt4+7tXmY71jPOtLQelbuDZNvZRkSWVk+O
0lgAwZ33BaDLAiV2WSqP4dDux7H4MOw9pjaHJEMmFo/PBAdWa7dJ0c/qhm6MmfRDCF5UovfkNEvq
CYTrhN+Aze3Om4y3OcjjjHUI8ZdFSX+P/Ndhjomfbxqn0eUXw0qbnrPLV1ijk4jA/QgzXk/XpGfz
+9PaICxM+Hx3DUsV+Ol/hMDX1jaa2Wwv3X5hAuo6tYsrVnX71hEMeDN/1yiGyCjCKageJ/afZb1X
ZQO6n+KPMIE83Tx/uwxF5REL3maeCC7MgWnI3doiSuAFdL7NQsM2y5qTyGscBnQzyAmwoUEhD4n4
j+AoqCmYNCQ1w919YUUWZhpml4yKNLvlxwmUfnM+Y2X9B7BqkM6DezrGuHEMlmt8alInQ8NUtcOH
oVvDdnWq/9ryWOSQsu9JGcXbKeHUOmMxn9fAz50dDiIwJHc+PXDu+toyvpr/b9j3oPZsuSe3Y57u
1Zp4i2YvNQGObgO2wPTezpcCsLNv6jZUvyLkHtpJBJKOmDM0TuA2giXHhxIW/79wotCxghgGqvij
YrxhHeulOgtUoQhfI8DCEM+r6yy7g9wh9bH4d6y3KqKqQxJdYa/3TcH2hAoGB0fWRk4KRCwxMwxD
JTq7yk/mUjpHX4lzzrkWmuLbaGoPyD/vuq88HaIytZeZ8ZdJ/VzWqm9z+ZyOpUw8yY69lFt6G3db
8rrV+uZuEnlTFowpE48eOkq8BVbhhWF/1UR/rAHiNrx3497tLRz5Q8dBSULyHHnh3Vu6ETxG8Itn
iOFzGbmhN5ahL7GkCVZafl3O6MAEbkPqJLoMXwg60iPDyVsDV6QgvmuZuRbNkpr5B5pKIPNVhhBv
Lh1kW3JsyfL46Py9EpFZtMjm6Bs4aBjgHk1uiitFcqBHu7hCuV+taALRVY6fqbW/DrqNvH1gJ9mV
7PQJPgcaWgPGXg6jL/gUFLyA6/7pV99MDNofASsC0TIpP8zMC7k6hmDudK+J22qchQo1wYygXQP7
//5J7f9Aem6CgBOWpf9U14qe3VCYFl3XoRyEMsTp8VaQMm1Ib10qWsAjChpt2Fm1lS1ZvBEznSxr
4X+AufhhuCEc4wnPJoq/vWHZhC0BlK6zoxVBvtBLB0nT3bClgKnA6vWfdS6i+kFKiKhFf8sv+QIa
CnZJ08pwy/Y6/kHHz9fQO4dMK4uhdGpjg/VQ8N3u945UPauh3TqnQjwTBPaQ3dm6JXlxXDc9l3nT
fx8POQiEJArPwmcKKuIBxcupXC+KNOk/7BgKEJ5ic3LD82im0RpaiPVngUimPeRXF12tao1arW/O
nTET9uP7m3QwbAWC1/B1msSOm2HoCEqLPZBXBTV+WGpRkkCpWjuBeW8JW7k/ypH/JsmMAeb9i6S9
GfrcTvT8cG4wuNIJkc/+3u+fXMjhhPd3pS/Bo2HmXc3jNNTc8fzP+Ho5z02a6KxiKlPZB4mUQKlX
ete4ugmTVV6f8f4H0UF4oA6b0Hglw9sVaJjv/Tm2w7EeTbc/N2Vbfo6wxAcK55DXVX6MC+uzFj1H
/gXz+K+10DfroDuiT5zaZ7yIM5z06SXrLX8QcfzDD9nzI4QAslTmhr2y0XD03UYjFEZcMCYQijJa
4P2nrRwMNb4I061d3sbF4h0D4GcrLaElNpiXr7QyKo+r9Hz6I4j3RQ4qmmP9O+Sa8HWv+nDWTNSj
PxdRMK48zpDtu0YTScHHl2ZIlAVrZDthM48K1Peuzlvw0+T4RKiz1Tc5BvEIdkrNrm5Tgbi+ziFw
PCUxSoft4iONGwUSYtSX0ZuVqEwbUPbYdyUaRA6cafQ+8x1CgkYBvRj1GrbzB/vTp8pBj7LjE16m
B4mB74TJnqTjJp0rBQ3JlMJUChPZ3ktWY6mL0b/AorFFk6m6HVHIsZ1pvkm2scmlOim59WaxP2u9
0tYegTY5ge1FQkPR42wriXXwEkWxg7rpBaPwHOWoiyhxIk7DPbl+FwVUHTw1E0OFTcUWtDznU0l+
w3uatduQw5/gUz5sL/fHkliZcyHHDrnIhmloseK+RkXQq4ROjzJC0AVufHYLmDvIe7MOsE0woiRW
AtGK1D4F/C0j+9bhSSr5PU45bojA/ylhgdSkuxcSs3c5F/oKckIO9ZXBKS/9hLKw+3RRGvxMd4YJ
evx6v44hGcII0FA6qrn/bYFG4GPgj2UF9Ll8RSDjCn8RuozkO+GMEL2GTwfmumu6jqxHq02eOXaZ
YPD0M1lOOIma6dCZhvZVit4LXLgRr4Agih1gpxA2uWRyFEddBV7Yf7fR7VOap1amYLdYSIGUPQIK
azR7v+c0JDUtxd85BS6SFy2PMHtot2X2W0foVDW+zrlcpDJyA0kPkQNBSIYLIUzX0Bjpm3JCjhGe
PYBYHL51nAhdGhWJzGlHbpn9+5wA63iLcMI8Nfskj31tkuIZauAKCxckFJTxbSBY/KhRBW8Y99rs
P+fS/zVXSjG2zT93EEU0vqoZdcrSL3hq8yZ8DrnvFFsjLxLpCDX8WVEz3rGGLjQPbE33u3VK163u
f0Fh/xIfqywgxyKkYKCQ1LIvpzDSVdXCGv+xxiJ12yYvd759fc4qcyvXF/w9InByCgRBv/+vyYYF
Ue4mOtyAjII0kG4RKyjMfUmwD5eGS9o/eNeE4XB+WjUtP/JBxpJS8sBYwPmY/p2sNkHuUGvWKK6S
NMvlGFs1N5Pve5vcHeIpGsTrBzqtUlxrNROjDMXVuPAhDQF3sfAu69OwthW8QfLcPbUpnR9j04aK
c6lKPSnZBfNcEpDFPfn5MdRa9RaFJSoi/cXHG0MqCYyQlWcfGlGT6RIIIMRhQ+PY86XqA/n2Ju29
XPXp+cjrJfxEqe8VYFvTjFHR8bWcz0UXItXrAQLfxdZ+ML8mBLBcKsqUSyrFZeTts/HM9opd2tlg
pX+PfhNIeoHtDqpE5I+t4vkvoLM1S1kFaY9eRQ0BX0Aj85uO5XYEYUcPAs9U3uEZhuOt/P3vwsLi
GSzOkzR3Qk3EG5hXGesDoV77h1ApWqo0aQ1p1/ImMRiy/esVsmN2D7mgYEtXzEhF/qmifqVnTPLE
MJFYIPXmQlBCqZkiIPYnk3vSfWqMUzr6eOOip04I+YIxVi8NLbciRmYejO5qvMuwX87GkxYQ9quv
0kqe4hqYCIBcW2JD/k0i9zrk3500nt/SJ27FwE3ZLVJj+h2saeM5qYWlxh/kumskG3BvZkumtUyi
Zzd6EkUINp8csep9UmjXKD8weWV/lsWHRD4DxvaTxk2El6Yntm1qjVO5hKGUiAt3vJ7HydXTyJCz
lfR0nBLLs3UdcdgXLMGXaExwAtTz9eLz9vFWzRwVkWTkrloLygp/LVMniHADlOo4+3kifVmLoeYQ
Sl9zot1gFrd1FFY+wMNIQKDQbjm4A0BrHm72yWGlaRzkmIZjJbiDV/1xXSpWtN/kJh36GNb0uRs3
tNTCJscJfb0B6PZoDr5K012dFNA1nqLLsL6hwaNjWq3rBdrRQlDe0Mnd6QzlD1l9PcdanpMyDFqb
BlOn3tzUKt4QOruI5WXFesWlUsIUo4V/y1lWxBBQc4soyOLOMJLukYOA19N9q2I3DwoDgbisshjD
AjDInH2kdL7KU/y7hmQPY9v4pm9VrrxFFIPGk4jo4khnG/2D49ej4xr90ROuTSiKSJj8kNyK6hzR
++cgP/NegsrHxXkR/Vjr76f8rIkMTu+cVJD9ZtUgTkMuYTCnrR5E3Svq1MSc5TT+H6XkBY4oEog7
Q382Jc/ILIW2k45NtaNv8u4ETJVZDsnUL/CM/YlUOJlqnJ5KTBkcS2l3Rl2TtpeuOa708EOYwDMu
rrs7n+l2de11z0HWlD5RVIPcZtlnh39Ut+n6W3a3NbJhM/fyT43Li2xNo2fM7e5XrSI2hG6V5wro
0tRIEbD9H7t2sgSLPF/tgtwyujRmh8DlvuL2i1z0wAnHhCSfDJBmeZmgpf9o2927PAJ5GKaC9ZuC
PRKv358xXFGUvzxVZdFhJNag0AxjJrcfO/5/SccHBTNrKsIpzJNTzX4fUwAK45LWM6kG4sDz6LRX
gacE4JPE5FDItuK/o68azKpJ7O7XzsR1Hky7okdgWu7AFy907IpfSTur3reevVc/XCYIREZ94MJD
dbqUD0Uz8A/uMtBhCN0i0ZZxsap/evnSEa5k3NDCC3SKxQxgMOkt/WcYsp/uLQTTHRYAlyYeOQy+
3s6Z8Xo87PuFG9w9dBGNJjhUkp49BcthlhpWsinO2YMck7n2qc7WkIbP1Txv+PI7GFTAZTw0GTkE
GbpU1VFxNhFu3BNdL8gYQZjwLQxWXx/hjQ5zibFzw3EYSCmbS4WZC+K+2JSja1gJcb8NwjPEAmOC
nwBFKDzdwTL81gpS2UD+lcyDyloI5U2xv3FfvWUqRX+HDIsSPFuad1irJSofa2m57WIjhZyobqEQ
oqC+hY0a4TilOisd/GbD7uySLlXNrorJjRcIr/OkSO45bFaJIusA5O4u2zq6mbg+7lT4JQvfFJ5f
JwHu8qme4tvJUowciEHVISI0ArjEm24Mzbyiomqponu+HEJ0CIqUkbxlC4S+aSqx+mNnHS2ixoFw
yCpMSbJV6V3h3Cuc+BnhRO/nMPPAXt/3Qy/KTpqJW+o3TKLUQPv34xLrrLMbFhYewiTAIZQBTiGj
JOpX8y2Mzjslqq6UxxoUvakyGdL4zq1lAvqjIfovVz9AzZCRvdxUDXDjJgb8uKNynQqVtrc+Jh6X
NA7LlpozjCCD8jbLDli197NDit2Y45Z3BjIlFIVy/dQ4yZSG4IgFVJB2sZYtEXGJz/UMLkoykASl
GcvU+WzMcIe7cz9HgK8EyrXjnKxXSqVEvOFW6b4ctymI5fAWdKgDpIYNiI2GxCJZTAAb8sVitpZl
6miQzV+305JSceHVyxIKSkVAQxR3b8KHRkyucAYiT0S7pMD3vqzVlUuLKjk+0Jkm06pOwbeqXc4c
glCfI22pZITq8A1pxeN4NMnTPEyR1tV2aQIoJ/0SQxioN876LtLe6V46Kh9kEnVXrYIrenhwNMtc
x2kqAT/WrzmISGcCZbeh5MpQpdDa2+KhH59zHiaujCb9jHXPE2DXQvKW1Atz07bfhXtYpVLfD2sj
zF1RngPL7S6E7CI+o2pzkghaKz/Ke6kz+xlDYU4wmvLkjYcfVCi3jrqbavaQXVMYyynig+EvhlEO
dqGaAuXK0SMfvVCVla4ccdkp5/cF9MwfW0SN4XLYkYUeE5RdcnlRwDQu/MLXkIkaT5YKFeGOwuuP
BzBtLk2csKdnZJiZxoxfdNmqJzgfJhyT39AeXR0D+8uc4DZ+z2mXPJRvSylWuQTiyEzonvjyT+AS
c5cX7Ih1KEXjiCrGGKAMvvBZSLldDkOfNHif6JXGk9JIoJtcyex2+I1WfZ3U8SIZH2jYC1vwMttF
oLMvCllu5kmMt/Sl9SA33VxCS25UBhMZc7ltwJLSHLl8jz6IPIN7lnWJUK/4x6ikEZx72SiI+cib
g7lOw974cMrpgRs8AwvFGSDPPpwwCPenLVabXi6Ty9ckIXZtLpsPM5mjPYUmax7vzxkbZaXlFlKU
qVxUtKqZaK8CfGSJ7CGFG++gbwQE1AirjtSmSetYvtpEiNcbmOujpe6+eNlYBuDLFz5dt7Wi2y7U
LqQZP25PuBq3GWT34/pflMmWTAfmVBSqqeIhENy4neFNnZMcJzn4Z27oaguKf5hA/YVD3GtO4fiM
8DFMgV3tvqCzDkmHWqqrAxF1STInWSnlHPAazjf2P8HZYpaJSToeEO+vvh/6NnFqYmTW4AaDEhBM
kYcShFJae1eclXZHhVs98SV00ZMGHWKgVW2tduci85iyO9/8yPO0BYyOwQezgUkUzCUBZ3O8tpM6
16fUgRnzd0zDhI/4dcGA8F88EJIrr+EhzPS7+n49IpX9T71+qXum1NRjuNuQkoNyjuAcVKktHx8o
LaNj2mD+u4d3LofDulKyT9ZmM13zL6BdHhhNimQF+YXKstoIuhxWvvKypYzb4FvPlSvbdjZVZH15
Tv1v34WPnKWA81E7VTCmIsc26ZyeiH/xqHHFa+mPiZ9RxAGzhbRmdhkX1u5ren27pHzzmb4BXFWL
zj+cHwSSMYyKpiL7UXf/moD+rUmDNxcHl0vQLmzwNeK59PhTPUqk3x1DuT6wiTFvfAo5lyYoLN3s
k1RVE8kf3CzVH9uTEQEFbd7qRNInJOLSa8ZU0UqKcOJRnt7MZYo0kaycn8cOiCsyX6RsGY6PNAYR
JXzQ9J35TGDcf/Ri2T0fuikVJAFSFeeNsIR+jHVeKmfXtswrDp72twHHKHNO8bdrSGPBoMxwUKvQ
nw6dgHmDgFyqsKsNbWUdan05wRXxAFlLsLMk4oXXv03q+rZJd/miHARZWNyG/fB20cEWtcfpJ6Pu
4IClIp3Zjj41iI1y1lN/CyEQzOZLkCRdMOZWTj0w/8EX6ddvFgTMocPX05DsMgalroOeRWttzjKP
pZG31s88vaLCglwJEaUKhalLGNNZ3OK87CGg+Foz6hIOhMcUiZ0hY2E3fxKsQUHxVP3t6d9CViDW
n3pEObZOusq2i8djMgRRaw/cU4TNc6OStO7GrzDRkn0xOm7YpesWE49FgvPNdoup+VQkwubXIrm7
SGwuadtpINwMPKcdepzqs1jhlzEy/Fyl5K/+/TGIjrcKhj89j4L3bU6Sd+jlSKNPFUiFf+oDrXLe
LqHSlY+zLggtygc5L6LRIU7f7y18jux0h19nJ3H6evtpREpZ/2AjARU1HV05JLiDpO9yXWKFhsk8
MSJhlM3RUCa8qCkP2LdDS0ODDhsdTMDUg9khWHOhRG6WcN8UgHVjWsKO4TEEsfkeNBqYkerlOOPF
yuLwqJnpmG/njLTPrROjadzY86zv/yaNGrehSRS+YbtvV8SQMQjMA2wtvhNWH5k3pV+S9u8m+3DJ
4NPJ9Ij9uRJcZty4XtWlFFOnh/KO1SOujkEKIh5vGktMRVnz6X4fcEq4uMSPKrrgd2chvn+MViNC
UvY5ca8ZI8hecWPV6EbtzMyrXQgNeVL5lINl4cZ+M/ZUCyJf7lhzWW8arNDxs+HeT1fTjEPJUcJr
SGN+SOki5H243jLh+JLudFxUtV7Us8zBajB1UrWQDQjjrBqt7w6agCsIprCj4Ovu8LKzFWFiCdXP
NOO5l7gc9WqnLoAqL+HiUrcBGiVPdaExw9dkQGryDgM8hAPJoQ9VN8Jf9C9jHvsMId2/RunJZuTY
s+60ohxqnHKZAV6wYrWuOHHD5pXUZKAk07PWNsAzd6mf6C93YenzvD/YmuiCmTaF5PSqIuKdsOaW
dE9DsHCuIUJTf4OOt56fvHDF/B+j8ace5+UMhl7y1gFsXeqtKgd5fzU1Svh0VMoTAAUbRyqO0G7j
F3QJFWO6qsoiBVVO+36Z5l5mUPz9oUUrAM3Q/HlmPbq31MCYomZ3++BQGP0OKy/2SuP2r6ZYkNm3
p5U9Cn5I2m/Kkt8O9syXPmTgFzau3dBr3dyaAc/g+KQcMPJ6VdLjMwejJipEmwnAaixEQXZYSUm7
8eMrtoa0axMw3d8BGUZl8I3jsNsfreVEr3mdJw4UKSvztqyFg+2c28bjHE9yl0JXxwzg/UfXVBQ0
Fs8zWq9yFbWfW4kpGmBIt56ikRmaDu74d4Ub0LghjM3F2AdFAbwKMpCmz4TPl2fWyEDRxy5M8Pm4
HCED2lv3Juf94VTC8CHEtHodKwoLEBSRDTwMF7SJuQQdNDr9C5LF1qQCGRNZ2f/cgVJHY0qNYl/4
Ad2HRfnlRJUTgLhHWXKw7RHX+y7UeOEo579ot2C31sZKDvpeef8FAEhs+MgY9+Hqu7TZUH4bmgfG
LDxR9MJ2PUPHux9azO6S1W79UdPX3a67b6cHGrt3wnWj+hHsOOfLQ+rxIuqV7vLLrTbmaNGJgNFE
4SZzPv43HrjG25FG/AAriTPm9oDpQPHnwfNhV6snAupDwfUDOOD3jzQZ3U15HUDexkeq6KUys600
D5YKwhaNAucXnvb6d3TciTPCh/qKeCpqPhbMDJ2x4mYeZ7LLMhNkaLBUhS4uXf9EiOdfB4Wc/doh
NmMvD1XPoSCz6NtF/8CixYjekeTZfvnCqBCY7HJ+rI3y3DlJLu5czSA8eO3x2Ls21H4NQtHTrgnG
TVTd2AxEhjRtcVD1JCjGKEzzPa9V8MGPlBvQj+IetAl8MuOH1cNBbgvZqtERW37yASTlUedTuZ27
SnuxsfAVCvLrMTyRrXOJHx4zi0G/wwczrrtlSrd76FgbedccsAsnRmYHFZphyfdff9PH7r5Az5OA
evXpVVhoeDL+jbn9STDVJtKUtbZgWE2m0trnk5/7V0phuolxrrWl/Hx8jBhjM4H6Yo1NTws1Zn+b
chedvd05g0BGgXRDYPrsavnpY3t1etqG08LoDhhr0SZvw3PjL9hr5MXgendyWcDGm3mbr9/BUwRn
+wbIumK0Zgx3OmkwSoLE79m+OLTP1S1YW0iRR9fyjCY6svVrBoUxd7CreIWGF1y4s9xO3D6jDNrI
/5UIUdROWBiwHbLBz1ZFvTIEZJuecGyDT6jRZJDh7A2bktNS5GWA2BtCagZHfG9DRKmEUer8vM/J
0krFBVR5r5E1/hf5KGBpxnZA/g0Nroheyu3veJSqgld+5y1lhckVkxd/JrobbGExGB1WoIWj2iAD
tEeKOzL4FqKCmK5NLPeZ9j4PzK3T5G+kKtry9KUTEhcit2ueJY++QIsvM+9RfeERbgur95Ki3Vmj
ptTwPgos/cSn3y+DuwW16tN93NCBs+D5hoHdZn75uHVv/cA0yMKgPkJZjAEhjmq+u8kQTolnGfCX
oafDtN68d5nwINRKbt0AE09HqD9sVSCjoygJzOKJElHXaqm7gFumF0KinhpTokYpGhTsA3c6jgRu
xMo8xFSwlOM/27qGZquXKX4agwbSRYS5FVY0z2pxgDAEG7ZFZ8czt7UMnyPYFWwJ1o8jSDhfjsEn
C8xz7hNplidhLfcjgpub38u5WohjmaTgQzE0ezZZIbHnznxWSWaz8Yo94juLaz42CuJPDV2RT+tO
uCMy4MtGNnw7nRPr+FRU5CUvQSnxx16N4MgGAKD7s7jXmOmvK0xOZUrc+nrfN36iJleCWVjLdNDP
Gf4jXidzNSQR8pLI4CUrm3F6lNy84Idl9n26sOko2n5/CMclnl/SFvZNoUaBfF3sUxqgk8haAqf2
dEyPDObi57NHTCwERGw5lX8WBfpKCCIa3D8G7sYWOn973mvVgjZeOJu0NLLlpiGXdCCkm8EJJFKh
llmIInOo0bTxkn7XeYlzu967EtUw6wKXenzNknw2QABp5p8iXjdvyEs7ylCGajTvYn4vDcixyGwX
9ieAuXupFmY/KP0PkeWpztOWYNjdDM3IJqlvTAo0D1w9/oUOqYQwum2aFB2S2ffJre4RqOzOfrBV
sJNN9uuW9aRhk0i4hy1NE0gSc+Df+Nc+ucKon3Q9v1WhFX7FRsxpZymyhMCPJ1mUKiulUo1jFoyc
1plsrE6fRTWjB90SakZFRn1CvNS3dWc++p6bEWhF8sFq1uT1Ipa+h5c41Qx4VRFrRggnViv1RB2p
YCl4Rls38d2BLsJ1iwbJXhRB7rcWISnMiG12F6k2qm6EPoF/S2Mgv6uzaDLQ3Ic8fZH77o2UzgSO
CY1M5ppTeOxCRraR9IWsg657dcCfSUV2aLLSDHeMs+5S6nzvqQKOOjCyT9RfVhmqBmWuyiIxtfUs
lNL/mFoYZNV+Xa3dOLXkMLKdHt4b+HnQBlqOPRzXqZnsuzxtTPm/vSewBZpBTmfTd3ELRq+V6flb
raq2LqUhhCxyijX25JqINUKJK+NX6IkiPJ/1+P6CpnyJR0D+ZQdURJKjiDAG87LbsGMZD5oKRfw4
VRR+whUTXztvnZybA83AMkfaK7iV0U0O3gu3FpO5ZbWuIrzJ/vDwYcMqix6FyB05eMEUo5l+eUBx
Ic3JMt6R3XAVqb5LWl24CwQghwttSZttaO+crB9lic74wr8k69o47o4TGa/yd93pibOMLqNg3Tvx
IL6xZwG1UWL+OuQhwDEzcvaLZ/WzTbFHXjEzNYXNTteMlnWKGGJOtFFoSur35kHWqpZervbZyyYU
+bbn8CIaHJog8ZtqC8cO2x6sFHXD/FMcKEy6OLVVwqnXs93hdEKYONFVFJjUL3KtVed8ZuCtTX+L
7opIsGnnbeMuzxM4KVdm2oR8FHDLnaognm5+GrbgiELCWyreTx8zI5iavpu7Fy929BWKda3G2ur0
G2Hkp8oM2uvIhPJLQhfC17dwF1kluFnofhYDYjFoIzgnmNMhl3mFB3DHJW1P4Jr0RqkTQH3LJDds
3lGiSC5uFxYbKDed0iVsx105HTcGPLcp8nhQzPohLZWE1wF4IMb1b6+PZlrBF1+DePeRTWWLN/qv
c3LwnGa2ZlQxZR6bcaTDIDeK+RkssMWRFG8bppd0I1fIGcLbFY1CP9xXhmrhgeRI3JTrOqbr2jr6
VR9TGix9UcvG3QYyHLSV5Tte3wYXgUjENZVtsZ+7hz7n9curwthy+JXypfq3FtAdzrm8ePGVovYo
AUwrwRp6KQD75XhD+/TgUGv8xFFD8LxddZZk70RZN8oJgscFfFYl3jEMZy+t/wMHLg71wEwUccRd
Sv4kcco7teS0UiyudXtO4x0RLDGZEEYIV/fZnPUSdRRRUqxiuJL6WvgqFHv/IU3zQGR7K5ghG/S8
zu92/lnTaJovwkkrRmoamiS5sOQXmeRLVGO16KzIJO9ZRkUROSkCD8A1NkFxyvrPldVh4aD4Pv68
Nk99faB4sl2BJudq+TC8/w/rkxP40rs5u15EHHCOGIZZ30kjZHwraOiNLC4cSzSA78DqlCOqkE1L
UhG+5c+qbBjeC/7LED+vDB0FsN2piRyqY3WkeFl/H4ll/2NwTAHuxKMmEs+mn/6xC4HF5Q0SrPi3
hNnAxhHe7qAFqozzPqVd9VgjKA0IEq/BJX+Ml80BFBuOcBWCK20nPXUV5uPZSd4qEseBTauR6CHx
7OIQVwZIOT37HLqIBVsbJr5Mi1mkYfsYIeypObAbE6o+h1BN9yYNgyeXnUSoV8pTmJVXeQAzpg4U
R7bDW+4c9EFLD+RJ4UYtlrD+NmNBaoBqzhmHQ67urtrH5cGYX5pARU30AcJPaZP3KjMJpZDf7NQk
1fVsVCmaJsfMPHSsGGolPAREzYpQOyPOo2FOsY0wh9QoW7yPqTdteARPGb2hSMoQ5iqaaeCby9Rc
QHHVKoQ98F/3LsLZ4+/p1/iE6RJokp/AU9haJqXd/906AmKEKdOW2mRNE6VWjjmeZBn7hySjO5wK
z4KL8+kwH7IwBEPNwQpP7TcIfsz0EdYxedIkPjtGYy5LiOx9wXxbc/Scc8kxXxaH5LvHTF5KqpEN
eh0WnTgBxTto8zR2KYtLcAL/ROxTMCn/WYcP/gEpZ6fMIBFzu6A8NI2bpP5y9NpANWHaMpeGNcrC
BxYi9XKC90heiLiWLaml+VF4EbJ6zZ1OtjIXtnXQ3j3q76bgrigXHPnnPlHSZSFejJ+LQWn6IevL
HUHcbnQM65BYX7RvLPU4iAgRNKMaffGuSjwNOFXoZn28ThzWVDbBaAKOxh0p+15Q+7cK/s87X5L8
3O0bwUyoVUv5yqqDj0AESpKhbQeN9xK6/wxzI9XmxaVaGIqf6HjOIkPhPQOAUfjcIyIH2Oz83xxJ
1IDY/F5ZJHv/W0J88x4nEbIGjNMUIHJcvaZBEEzEOkblq+BEEZAgjvpqqb1fe+4U2fYfCRb4UQ3x
EnjLunJ5KuBEApkdh+sMbeluvzNr3CLBGEFgQEcztc1KzJyaAe3RR2RO2VzWU5EOBxcwojLrnQ9d
hr338jj9K5aDIdkRcoTRs3sCIZUgEn+ldVJYmcZFNaBAmf5PZg3cHUVeJu3RuQJcfw7/wF5SzbLU
ssVeMDPeSZxeLP2jbjHgvvK0PWO5YCCGWrZON7IchSEZMuPaTdqmujPL/3F/Q7DEHarx7tJkiGMc
Ke9EWrtyhv9t4TzgqLdemOW+UqXKZoTItOJkMQ7UhUNZAtM7CvRWPdo+swL8VaK5cS+cj/JXlQ74
9cmFRzFnng0tjCHEcpGCKjVJLQy64FL5aWTjc6UFsNn9lgtbn0A0yxfTUGF2jH6R7ygjPA5RW67b
n/e75V7WtEoNBmtbr5JCam5jDG9J6RvB9xx4Xo7Npeu+KYb0Dsh9jyTrreJdD+vODihSu0MmyYnD
JOUqDadbkdozTGp9HE+oOUSp2V+G/aie3BUj9tbetLIJDQUWQlq+Psp/xyu70ESCx5vmV7DMAskX
tRMPGgkvb9+c0iWyZw3q5ha5Tc2pxBbRgmE14/96TstKNF3FDxZOUzDqq0H1Fh1WCPpR8cKH/QiY
c235JXnAPsffo6ya7z17WtPzUCfUkY5ALyYKs/L5F80DDex29YaM9shGtn1KBxxfNt0yxVusphJ6
hdIi/YwGd1QUiPG7Bm3hnu3s0/79DZrUJxHp6h83St4zHRekaAI/1+VEd5RlEISDvZlOM0fXueiF
M3eQjlmMhig4eOwfhWaCVel0yotALnzhgaZGBnTugvTdwt98jgmUVojcRwZlkJ1DBlpTHrNAb3qm
k3bN5xFd3THNZx9rn7TGxCsq0AAPl4W0GE9oZaLRAtL6fQWHuplr5bKuYav/Va2nFNazDtUxOjpU
tzZuCm0nZI/sZIa6RDScyC2p3bZAYodWyzmDhw+GgFbbB84A+4iwiCBdEKjyxzQ6Tf+adD8WBn/X
/gxF/N+dEFsVc6MzjKOXtEg34SN/KS4YDkDbAyM0Z9HZ5tX9xi898ZXpTBJP5rxmtWvR5Il5/LYb
Mah/Tu2Rp0P6mXJ21bJm/GyoTLEVLZS7lm2p62PUrvXs1Wbf9zagYoCL+FJWtTqqQZhtCQHSICiz
JRbG17AdCEc/QV6NOgpZijy96jnk0ms8CTK4jOePsDBdKS1su9fjNy6SLdP0ZDDUXCnwQKojaxkp
4TjRZyWY65lRSxx7LpVfNYmIErDiovsJpWqEEKVXdw6dLqVUCJJJ93awfaJG+Spq3E1Sz5/j8KBq
JsuuhpEuZUw6yzMy/xBuKogViX0zdExR4DAZFB000cONusSH1hxNm4SDroXOdgCwUmNKAXIbkEoQ
jdBGvFelI9avqqYoA7B+SQGeTGZagN8JzZdfS2QTyqpNiZDQQXrlSzCVse9Ag2Q867Y/OPKrU9dU
hFCkP1Dy2skKIvUrqvZGavbNQUKxkfXW7fKNHn/hNZJq+ueSUJ/VtnnhpsvUU/WXhV1Ifu0JcH5B
6y1v5CgTbg8RbE5iRnK3Q/Cr0tOtwbmjG+tAimyGB5HImP0zOtWr1qKM2ndT/NzjgPLg+e02zLDr
PDlSaD0SAYOOIM/PBiLrxhMwCTqeT71p0IWH+mxDySWU5r3ggXa3tOjwEClNKccbUd0rHqb/CNHj
+QZd5XITkjs+D96j+KrL0WMNOFwPeAR0y4pNuB4puGzvnY37mpd7tgfI893PuGbbI6xs4/ID2UBY
Q9MEf3afr5T55JRCYuQrBvF88y3oREenNRX/rD+vV7GmsDHFikR+uBejezhajll9lKwq4oEVNLYc
oSHKtf/i7jnDCSEVjXCgj/hg5faxTITI6cDLEJjceqGez5KswjwmNI5w3h3p0eNF+qwzblg8qaVe
uMojk9MyRd68cRK278g6nohYcMa3DZxnakU1L/+80TqZjIeQF7XGqe8WdNJblLr7FxgydrUgLrB/
xxfFiZHPEDi8T8u3610i5THqTQDeTggn5SzoQzYmAYYl7ZtKcQ8bUu64SArwPvGmGZ/NFzrQTp3h
A4sK8e/3zK5fsPhDN91tIqpZq7Zk2AnR5rk03/iI7KluN6lMj9mAJhtldXlSHDmYqmm/stdVnTYc
yc5dsX0unAEEMs5WZu/2UuWQ+6I8GMFzSB5ZvUcRBV2w/z5KSJHO/5hQNIpByxrJjn34PC492VtE
vNOJw4dnfvwP07vgWwX9Z9A0NfPn+L5frG+TKIfea5As6BeH0CThJoKoBckCpuZr/altUk0bkGMP
FTPNzgTqaFnpuiibb7qZzaPTgloMPYcR0P8qgD5TgPKX7HZM7iB07+mL7KsQV6bM7RWqmk7MexD5
yYTHHJP50L00BJM3KRlfomk3mf/pZTliYW0rfKRGxMzxP9EymXWrL/WVnLDF+lhqiFN8dnQ7dHT6
AT0LY7IMhAs1aAZ+2G2wDtIDAkhrdP9J9aaiS1r7Dq9dvVr+Zwz6Yf4rQmrOvuPIcjvWjbgUGE5m
5uD9Oo/sJ+FcpvMcdD3iqcrwtTWBgAHZe4Vsl4utKWqREJO5pK42ODkXAuM4u43E1oYQUNWjpzos
bRKPU9PCbAukFRCHfo2YAtNFxwrwQVu+78xd9cfAzUJbHy7Hk/V0U5ZqPX75WjSCZxXHF0IP6ZtC
A7YM9U3lOVsM6mj2IASxSyKOKlHOMmOwrNeC4wPeLSUtRErgacdXPTomnSbcTP7tyWCetdetGk2U
FU3EpWSCll6ztaaEDBIlHJe8y4rPQVppwRHTaQ6KgS7LHZNdkwxbhslmGDFjOdGGNO1MhSi5uQkf
kqCnO8zCrdQ3jCWVCVKBucqIgiLnEn8Q/48RjaxbxPjFo5MDk8BTqe3L1LqRLCaDvzP4oczZqf4E
NR/x387EsPUNIbMusf4mRmBhtuoDp40J4KKm3LAwfoS/tN6CQJeFEg+15jIHHcNoQ5Zf52Mzac1x
TTSez7CKDn5dKd6MIUvqVMxQ5MKnnM5QSqUQkdNvmQjCepNDhuJCynaXszkK8C101ZxL6kF1ppT7
+4H6L3p7pT2bgZIKorTb6iZIuI2SLiE9g2i24+SoamLj6qrl+kMGeoCugf+t1wRAjvuCqzyjbyN/
j9y0upezUqd/TmjZbncWjBU/sKsfOFkneUzxzzlJX6X5tX7Ihw/PFWQqW2daURGZDOu3OloketZo
Q6X9snLK1PZzEGQrVKktbDADq4wbGeia0Qa9A2igR/biOq8QT7/EH0OkD8tkVG8DET1lwvTCpQNX
vZ53Xa8bnKCijcAywUTYfUPcVTwSrn1TRanKJosPtAGztZ+n6Bv2e5jA4voYW0uGWvpkWzpohEEH
xP87JDLe+Ynm/0JAOtJi4pt6M9CYkIQH+CWo8h0xmcYztUJQiwxXMnh5WJUpJadWqnggvpcrrGQJ
mxV9zC6+OlT44dzZjHxFrUcCUHF0hiNFrqi+WDnJBasbeGDUqVR7HJABy9IvVblp7IU2UT0xj4gj
9mmQzJ3IpjP2lfQXnZ1nuLWQamEnerq/W0LmquHjbJm/G1BzF1g5fVrYSJRmoQQHKDEQ/Yq4DMI7
u0yTGqhkb55VmRGGrPXXNgjkjeg8pZTjrCJLlQqca5WoXiL8g+y7b9/giUX1X0GuwfaWLmUpjoig
gNu4/Qwe+bJr0ZNSC8ACWaG2Lso3w4J/ht+V3mff7yAE6UG06apWfuqVP0LS6dOnpjq8PXRJMmDq
U3vYi4GtcigU5vWdatktPpIT9MWKEiZ+NsaneDTLfkUFWWBfDCIreln1lXs3LEEAFwFhey5pPSwi
QCXqATEngwCX8a3PUqg22Btouofs37E1epqydqp9Yk/rwoK/gMRp9/nqIHF4ieU3MkUibDwvJU+B
ASEJ70ZvpVvWVDXA+P8onGlTj51j7VNQLW3iFOXxqJ1mI4Ve4Vd3kea4nzmR9CN0O4RKpQIu0QMa
C02IHJ4MZA780sZdJdBtK6Lng5abTkgyFe7AuN7XNEdG/i7bCLws91O9dPHV5ACu5wBD1dGppZyJ
/fJwxvn4CSIepH97setbW9MsB5Tnf7XVzk77g0WC4vfeTA0CIfc6+GzXBHZ+GWkWOiHPw7nnWj2U
zcusLcHlmrQYAi2WjWrtgGL6ptkTQEq7ZxldAavvmOr2ker1Er+ZDWj6krKTG0+vh2h+1rVzoD08
gtb8sqUXmImpcKvuZgkpIGLdIELUzj9A1HuGd3g4lU/lWw7ROK+4T76RRPrXhViF1QaxwneHPWkf
vKBQAZhBfPrzxrGfYsHWamPlSqKRzjHD1JrSb2y0khrSrLGxm/SdM+5m8chlb9vEcGNmVU2mCIQj
2DwszuAndnsQnDJm4t0IDEkuE00fepb3P/aqMzgGjdS2z+7MbB8STwTAEuj9TMW9qZv02kXHI7u1
ndPan83j9Wjsfc3v49EUr/klMnfKiZCDSFNjd37fpvgR7zUrbdnd2T55GFALA+d9pYmjfYRdnmuF
lZY/gfkJN4O/cDGL++0WAl9IVCMIsLQH74DMudezMtv511VnuYZG2aWrIjTF363NZyzPLyGvqs7G
uQLa6+H0A3zY9HCVnfL6mvXihA6H70oimuAST8umwWpirzc+ZZg9JX7maxyDwvoyKx77g1WYYAQe
HAjcRpZbxXcS3N3FfsKF9xOYPzq2h+ZnH+Juu85wPYpomU8rXpZp0aPYMnaY39sgVt58wR/QVOcu
h0IE2B7MCrjkgG5vQ5EuEWxgVXBXxXrRqF2TbvIKCUdnwoEU+0bPpvV/+OsyipyOGu+klukvXh5c
Bm4GAjEGcR5Z24T77VuAM/HxWTmXHMHjwy7mN8r00D2d5gm+AhV4Gn1K1YbRRPFrPSYEQgmGjJ5L
hCkG+rgLdQOHEPTtdKLp/rc7xTzdUn5D5pERztZqAiveVe/nQCp62+odRtGydD2LxshWfuvkzzgn
5wCcKW+CewXYPPNN3cWVRXOs1hpIpPero0VBZAVxwMfqd5jY8ICJ8joRxYwtHAqWqTWbTLdcuH3Z
8p/+CyAO2pE2WnS4PkrQ7kC7No7/6UVpVsHhF8LIjsJuxjVQEi7QqhnD6mmwqwRErIua7bMty6T9
BlhsH390bnRn49vxoo5vNCEfyQIZ1AhZNaw9RwAHQJqP3YOe3ySJvkK04W9MLJoWhBO8F2Urerd3
5y3+CpFU+J8aTT4clWwyKkm4DnJ3r2x9/YZoaBgkRD2GInCkm9JJtgJWqYyu7PuaBNzdyY6Ivn5f
+mtruCNdr9nueR/FOlQkqS/sP0FeEWxXynw2bbePaXq2sX0VdxwaTkDxnokjjGJ3MHuwngkYwk1g
vtFiiWexc4tKPf7cwnZzL/MbNvZ6hpy0uCZVHWXQJK8se95AsptL4XoTgWE18YguuYJBMdjdRbYx
k1B4kGF7MTqOJomgfmJX0TSXUy1Wq5KR3Y3EQWy6IyfwxHNjg+0X1Ml7Q0jsyVKiNRp3QOT/MvJl
TigNCYVZ0Ln6nQSpaLpoN+BXde2NYws3aVUU1c/twuhHSFLMAHOsNU7aM0v02cTxnYBvaKXsFXrx
zAhtWYLdCWGCKh55tY4h1T/V/irOhusFb0dwgP8mg40H2cv/styu154f7599HwC0jTSHAFUua3ZT
to+pnDFNAoGOnrYYDJtlPf2U/layAVESLDCt5SuB88pyTp6MeK7Dx+3jmqnzYvOkSdF6a4JoxTkL
AOKZUHXafooVCob4+VsYFwk3hZ04oDb+qg90N4CA8OSIrW1icSdGK3Cm2Wd+ldmq7Ef3UCHLv9Nn
O5eAEupcQquK5iUSLJx5QFMqlMbPcz2aRa+OYrraAcGTzJ19Y0ud6VTebtWjUhWwshRJXvQThmSk
C/mFIcSnNRLaKHjfQrECJON9FALrqh49U16clkyP9Hcm9JsZbEM/gQtNqsG3XQYlyGMObO28A6xr
6CMF2VkFyc6Tq3A/AqIY8yzJLk1m0FUZNeDYk75d59hAQlVxkPyqxRYoqJ5T6gjWXgeWVdpJB72Q
lcaFohwBZEVWprIM0heRvh/jVRbCkk63EarN0uNZ/d16a/yc/c1LBYq1h8mvuw6gqUq7JIH9z06n
LISrz9FsT6EZ3E0Ur/fDxGQuVBpklc+pIFRIDw7GnvXqrdd2Kj/RNWJtMS2Xl0vGM7Te7/QKRMS3
jI4x/ZUqlA39BytAjRuPIBSxzaHtzhzrMsIbCHVkJSQ2nM5stEqIVAhvhjR4kgovzpYRkquUCUUN
zQa057a+8AVjthIJux0Qc0C2aTq4w0OuOU82SV9R6B0Zyx/vpHZ3xULUz6Dixs38FtNeOe9sth2z
qWb363DHiH47BX/nEDzQPmwUQTSAlvoDkN0+LaZtJg6l6EypyBmZYSn8SwCjcUk2j/k4dAXOJQYr
OrXEFwJnHb+Sq8HHrXIAFTwyhlD7mcdPjnwpfrEDTj8opEOYKaIf+roQi+JcLPvi1MODgN3Mb8FI
iElkoi05B2gNKeh6+wOggUSxzBoXODa9PP0aQDkDQHB3h/irdM4sO1bgKy7vvU4neybl5MxA20JD
d2lfzEyR+W48FBrIQardgYjg0eIfzmJYvZkDWJGo7p9Es2i+0GZDEl+suETeMyu7RSXVGWKrG0DK
7kqBuffcHfBHexGnOgiWVoYz48re8Zymen6Hy+0lh3OcNImFh6VwDkfVIP/xJVauFSmY+0jCFbmx
+F9V77mMlzY2ZpXqRr1TwuFWwJNiVAL+5BEi+wwQ7L1N8/IOjcJ7ytAb/RUOs+D4ySkn5feHDN5B
ByVQpUg6nIKaE9CsjvkBtUbSSO1kyP6Z9s49nX6Tvm+B7vp/OcyccP5h6pdCUioBqYX3UnDFKf06
BOYwm5uXaZXXY7ZpJi9YaINg7Jtx0lv2s4L6q+DkYCnTjcuoyWot2DpgT7E9CSk3n2SgeAzuyzAx
bq5bK2JTN04XS+0OhuUmHs6wyDzAGjC04ipjNi4UilUAn70G2b9JGmM/PHbJuSPURexD5fjJ6Rg/
v3Hn1AO9B5zNnH7VYqEnPMTvyEMQ7dQIF6KWhdm74soOaeaDMLDklpL8/jfh1u/yND1yVmHJxPiA
IivRLcMz9cSNparFncmHbW7x0WHQWBZQrT9F3NlLh3bOvSbBpEbFpS/8JmDd7QEH0t+wGVsVNaew
0C25nbZEQP5EnZzHr3zvZwF0Fs3aF6p+do6A+OmdULq5mWrNA2KWt9XeRMOqI7jpzNoE8BKyrG7S
XluwZh0aederyGkg4M0TYyV5kDdIyOqAasrgXKud0McjEIpc0O6tcd5ANx+g0Wolz13xYomCtdiw
zyNvudGdDYS2X30rRQu69OMoZqSjLUQABG6aZELfsedwu9KKDCJNO5HCurvt8MWUpFEEcxNAIaek
VzkX7rdQtNCAGdbQud4ZNNW146oprfpT3gGB1g9yfXkfMgrgRXCcW6C8K/u6+yfX3+zR0R8oFZBw
H4YR/ORuWyteGAk36SHb0qhOnutvSBgA988w7Fsc99yLOngKiQOrxIZ/E8JHWKt3UitG+dYZm/5T
+/0LvzMz93+poWWB58jR8CWdcoiEYqVcTQTs49K/cY3UQK4CY3xzWLFs5W2TVFj6LrNiSHugGjGY
hsBZeTwq3vWJLXMXwgwGfpLtidYLP2BL8XqBDEsrKAXbfHaKRWOo+XaKuq0Jimu6Oer1BmV42Gy1
0Q0hOeNI+U2Xu8JVRWhTyvntueV2qqCifwxw7Sqblkn8PYN3xDSIIIys4L6glOLQmlK255NuLPgz
3dQl/qmOfJcV972Ds+1NE7aAhHNR5auSfC1MQPhTP074PYuYVISInZWt6vdzTmNXhy3D2bUt8TTF
8tYaxkeBIIyGUvXbaD8p1rsdjFJNYwhMg8Q4mJuMCf0l3lFSVtypereRjJJdmOZVdEnIRC8lW4lL
vOOWrIY1362hsppZK8PDBFQhAga4bl4nEatCyNHHPFPYbjaFffZmCZLH3Vtz6szc6w9SsRMqnezW
F5tLRA2K+qDeRo3JV78Efmch2Dyhl8uJTIbpe7RWm9cmBJ90Nt0GnJWDW8VbybpMa4iNa3FcQ39D
sZ/rwV9g1Bd7f8pJ+QNxA9oOOJIJf3dLvtzC2ltt9zwLr7xdxRLtp16+ME6nRoBx1XRouyi5UiTr
GmZTH8Fo9oa3+BXrLt2gcAvS0SKGiwjRX4yXdTcErxl5m0DdVlINKRr8JH1ve15feB+6BhxmCaya
oBC1sVBT4dAH3Y9QQFGDWyEUhn24/AcBIo+INTWwhz5jggEQXmOX7QdqzlfkDj0OhKPf+z2xdPNU
tpEJg8n/0fOsWsg7sV2L5X2n4IKNT3mem/zaNnoXCyxSu4UhPPbr/cUXOmbE5lRwsZXHmNMtEOlQ
dxMuwa8ZAMcpN1S6uU5OVFTWyAs4n9bWdcKMkXAuvhb1iqzuHTdGHJL32EZZcza9xhsUfduXvet6
FRFKpPwASOtr1AMktJrmMaqBEUiVwdBNy4SAWf1dSBzGr0/PpOujzwijXZL+pJ43WbR612v1z4Ai
02trqHcw7lM3ZkrALh34uaZ7LFiUoC5jasGxbGrB9Zh/OxliXGTNrDAo0ntZGDCgmbGzfshn78fl
HTtMr2CdTu4Yr7sSGL3JysDSowcaFo4Z3vo1QuPpfpRENgT6BhKdo2+MamWIHgUWgiDITsqwNwSd
I1On+UXOSQWmDc2kFegK9S6cM2D3ThiqVD4cVwuT3BwU0Bh80qJH5/IU4LAOhLMA01FqWDU3sTPe
LwNWarJ6uGbQuhLk5LPmLJJbFki/FXJVuntdfK4cEL7FXbhX9RD7Ns1c0JeuX+/wqIfLLgOehqmx
X1OUzz/uxfHt9CWaXNA/CDMNhItSp/DfzeFRiq/WGCEch3c8xfL0pOX8/uG6NifHT6vHicRrk/qK
sLYZSMd+ytSR37xw6ujOKI8FxcsQyV0JqjDEIzL1TPp9md9ptnce6vlgnHsBTShcvh7z3GoS20nv
R5TrD8InnCaw0VNSEvfmaFJ2jWkZDtzfO8zgVQey6zzBiwD0XZrhB5Bis92blon/BHmFXF8D/aHw
WlX33gJRApAaye0WLs34UC1jTj7aPO0XGVtlU6UUC+ce3uW+uQ9JQh+E3DP0qWdvh+nk5idheYP9
n/tzxlVwSYCpZGXnYYF9qXHHKH+/Sz0U8xMBL3wT3E5nF70OTJA/eC46uXU84hAjOS7E3TIcIifu
rOO71O37YnwMq3U4yKLsu9ZYvPH2q8J6SRozWDpSYe1YFS0J5VOmuYnnPtJU883rFCnPmrdQYi8F
0sK+CUCd6t3qY3PhIWm24k4c8TpkKl13nahzbcwfteVLWEurLoC38I1dv52l3ZZ3QwJmas7A21Bs
jAyd/Qv+byGzE5Kbyqlxcpv/pVE5jlqJRneMDyYjvlzkdUBD5Cq7NPaSJGiINYZNsZAYsdb1PSDy
xUAAuRxjXnDWDNw06e8GeAyZFJXSxdQ+yrIWB78mky3bAS8e27in84fikDZeorTlqTH5VPUu8xAE
drw0x6G8s+t9DsONT6X6XNHC6gka1FUctvNPuyDgw/RbaNVLe5ysU2IZiisP/dv1oGcgbeEb8HPD
THikUf9uY+RBN4gO4vfjycEP2bRN37PxPfwszH9yrzRysQ+IgExl4l0qvZCAmmg6o6ic+KbiWboG
MPgeTtfiuN8vcxMjSU6vaaDNn67ugNR7X6PJ7x14Xn1woxv5lHov+duB+CY2UVM5faELyHA2a2AN
z6JJxsg4hro4WIj+Iz0mLLGQ7qNVgX3VbdYybaVkW6jJtPNGeQEE9Li21SsZAvW+OwjOVUH3FniL
VY4c8BfYdCW7dvJXmO3wjPIHGOohaEbzxD7/q6vP4X80In/VzOniqYSkG3oje5zI+FkttrmW52YJ
P8OXossF7Ye28gvKQUBV7jtTvQw2agKyKPvz5hIDtz/J4v29McomscX4JfIE5FkMaXQBh/wRusd1
VdpEahQeUvtd/uTxx2XrBPV5zuzoDWd8u0vCUE33Xr7ptKenSAn13SZaEc/b64I8VE811InXWzSd
Pz/7jJkdbtrvCXVptRXD3+uz6IRc5lTwO2KFnxOaeUisJPSOFyHMyVpvykP1dAQsTUUg27tUrBD9
2PzAEZiboenXhhx5p9to/I8c6MZUFMNJRAqeVZ+CfmTruDa+DgKVpgg+9JCZ8yBAAsnG3ovUoR3s
9ikDESbt9LVkSoDs01lD5LMr4LUR8aV8nlgwwHkYrIkdT/CE5bJT1LySPvdFMfdzfJ2H47lk/aou
GRwz16M4QKC2TgPKXYMVWmeUvkVtno6o6oSrmEEeYWFD2l5dVdRxdJOSRDwsfCgK5oq2Ua41wiMq
kCehBcqUR3HRqgxOxBoudBhvJ0ATxXubjGe0xtU/fL0/Kby6TWEmldiFTMzScRXnrI5B6b/eCdVz
tW5xybcMJ6I8ghi8q+OWzwT4ZJlpeSTEUFyz84fKZKR6WyzpjYznTW5xcs7DVPybo58YADL1wH4U
69sMvWlor/+uTygStZd5aixN3Z0p2HIK9dQvEa53eMM6y8DSCsDsjWLs15LHHxbMeOhBsI7L6bxk
QT3+7ZT/1+4pKGXDrdbLSUMHuORC+yntiaj6fZYbWiirtXFMnUIvqUEZbjkv/ZHmWjXi8/KLbtoQ
Oi9yXZYZuzZ5aaDq6iV06MGJU88hrgB0DTolbJmcJ3Fx/bF9EQqCiflI9HjQ4tibtvk764RZM4/c
xCTdeRcVoCxykTlCQBbyBM+6Zo7razKSoVGyU3ND8lNn/qX/EyYBKcmbZAvRz6s/muU1HX527P5a
dlDzowZFo7WC7JPEdSARneaNXnZgTa79CZPzK5RPKDiqUtPvlN7EZqiG1H/PgzQiXCA61lDgHFI0
Q65bCA5sTlGupVO3rKXEHvVXfTkdnp72mieXG0hQ1boIdEQnRladD44Gtx26dqf9lYTdX1gHSLI3
xFHVCBye4abMCQoYO/jRmyH5Bvj2Gst49mrSMcbHQXtvC3yoSmUfxBvddNrgFgmqnbGsRBXyMRi1
Q2dgEJCS2uBR46wTDwex9Y5K3WJQTWWhq7KzKc9t4p0+Wi8Hi7DVG1dPw5MOCtIg1CYWELRy38q6
Qgh3pmIVgwOnS8t7HFG+D03pwCIWbqwxZoVQ89yTxUVgLknQ0eYFMZYzmo5lCgVmls+eyWTNnh6C
oeVRXAhlnQzE2y8IuADIiqkXVvwA7ndMdLLIuKHnNOHijpPSr0gVeL8zAOu5u36CjwWWsovIWtJr
4hI8nSsv3rrqY2ychg6DCI2SJZgidgNHwKJnyQLFWo3jKtNaCjelSUjn/Fi07rYdY5olLUIlccmx
qxiI+ilhthdo7ykmMxxYRhBsVqlDHPRFBixzMefp6d9pPpxYqm3u4u5RpnJhMUM8pl6fDVJShJ74
tmA54YzFsXWuYHNvD5k8f6rvbqUhWLsrgWqpEaKUUyT4AfcMMZyE7zzljmYjBnqzbbiicrx1Hq+l
RVqT0EL+JP8fzujAnY//a173H+3vjG8UykXVqoZgoQ4Yx3EU+1j50uDXWdEQDIAh8CCtYz+3SvkY
I8OZAE/UMIfTEBVayhnpX2dzAmIy1vMUloA886bm5oHZj6Z4DJbO11rVpLA0Ki0GwwcoUTlf2ng9
Ccm0x3IEuokDyxlQDr+3CoLqbhujg3xaWZjHfa49Yc66IUWtUbxzBrCG8lz1MfyD4M5/bIDCo+fy
pCMptqTUew3d+OzcIWMZi2/uTt+tXzJeARYZZ1Iyc8JGDvrbgnkphwuX+p96IBPpi9TZTbmWfwDW
eODym9NFN0vDb/gXg95KMXqYSAKNk2V90nWHGJNFWPjXvK9igFiX7VsxR5zVB+G9WYJBnnH01uaz
fKdxIROtQ8uX05kGStgyRVMxcFRCYYkhWtgbBJWVUqKCbNWk4gEq9gxZA6Pee9x88yuudvMVvyjh
x5YlUJSOMZiPW96VRWqtS1I22VC39R+eTuMi/KLi6CXSBCQrM8bULQveelEpp5CV/dDtEjmuXc31
SpQ1NqjD3ZbNhalQby+igqWPkJdb4yIMUDLoSE3/ciprWWFxOXGNHoC835s1E8PrtoIm9h/7HAqv
+RZwAOgoWkiCc9v8h239HlJSWh9ryqD/UOdq+Vrz6ggcmIpBWChrkem8BXZOEazwaKah9vAod0SB
HwMBmHXn4UROljDMPhDHtdSbqgdP8xx/nMKTwB2kd3UVMAgSwmMiIqDSpzbXYlpnl1kGRD/JsiLT
NPkHqHwYks2WVyeG/m/bB3HSSv3N7Ysh/y3i2Gi6ABr/COcclr1tOViMhaXslOEUarhca7KxKwjj
CTrzUgxOfJuLYqgIHiSiZTNBXqriOWSEpCA8ebgLr2YiBRxJcdrDa0/IjXjn3Ho5sHQTl9j3Z9sP
Lc4wkL6Rhh+7gM4FIZG79Yt0cjnSfHmeb7/Dz75vKESThPj5ffKhbwOJMRkyOaiMS/7b2gxVNg1o
qzghG/OhTwBzAhHycGz5Csf4OsJgaTsjxLRj3s0V/I403thHa/f62EtLdaMOL7s5fjMzPn63yh3v
JbEEMkDDl/C0kFBdLRzh0YDEH/E2onIzZYGeinOMQV9vKelSNd8in1pMwCc6sUCheFHMRhGZwcXM
m4GS+RiCvkC2/guz3giIIoSb2I46+Au39Kb0ETSxXzdhuQxjqD8AqNxwHK3oPXYRq7mP+C4ndi/D
cEMi9aQ8XPsh1n3/iANggCamg0JzxP92Vo4Yl7SgXRCOo76Sy6gtHaYwKISnbaEaa1SwXIiPqpEv
0829SuPBaePkdmaCBi2muuBRWG7u5EeqsesXPfxQcQLHQtoOsOwmKsdcU+Lqa+mUv/EEJ2n7/+Tl
bxjUxq42ALX4q3cidDFw+dofvSK7mMRH0VWOWmlBi9SNd91mlIlp7+gy007kPJ646YTJZsrJG5/E
2Vf4YjqePMJq8qPeF4Vv/W1Y1osfD0pkfhDcNGizaw1jNFqdXWR6ZOEflx2KbGq3o4oaPURx4WoU
qYxJhYddXzHZJVj2h/E00aQ8ez5QjaKnsSAAJc4YrjeyDcZyg3/LJlJ6Io47+tDTGcD5/VqtoOPz
zyoZiovUKIBhKM3ucnS+ol5WZczEKHedvNa6r0THL0oyr/4yKuu9iieOOHjigoB6rgEKWIDUQbOY
TnygQ6G5zTWo4FdH1wlsBhynLBuAixOWTrkfoyF008dGWt9Da2lwpRHDpgZddZtTNgpAebHA1pRW
CwzcDCGlToaaqCga1oRDTm1vCLU+oPHru0vlLwSIPBkooIYMxhCCyOLzLDJsz0ixribX6uviWWLw
qjELDGfLOK+LrMEJxjI4VKMeIfGxy0Y8A7lQmLAKNWaETZfH21bctLPWNCYcB4j5wV4Oei4n1MhK
mUD/kf842wDC1CeeWX/De4vk60x3oBhRzP8ACoqcy8OVLhC2oR9i8U7rGm0Efj1MI7xet3iWHD6p
scrQALjfLlRmcl6ABsgHt3lrckVSE2jv1heBvgKg/wAtUwF5uju3qCZdbT+A5aF6cpVzndyHV8I8
dQJtDJOYMmzOHmsKDm7setvHLpB3Yl7iEqGJuOHUtlnBRpRO7gNiVOiojJ7uKcc/eKyNpgeQljEB
8r+gi6A1Y537ge7/ockQ8I/g0dNDR3dw+WMDrM/ZY2rBL3E2F7ZIe+REUvGQDyJCe4oHNV1FLOZ7
X5Tc0vENghKZpZpPMZpTH70rEQHqfxc/jXHNE0foq3Z7N3CbCUAWuj074SPNee53As3ZZIZ6ZkcN
4UupxJBn+7xD37jkc1DqMACHAxdu2Vj/FXNfrkmJ2XoAX8tfvOX+9OQpmAL/rSoXzTuh/OhRt9IA
gbhI3z2vz+WsakSLmSFuNWZttB0+wvrKVQ/R1z6r7AlGcJzfVjyn4cKIMFBOSms+acNEpk+8tF3v
5qBUdxSn5phqpxsEv0F9FpQblhxq/mFto3zKul8q+1a/4WFpxVnICuQ0SclsJCYvbtFYPI40VFKs
lMVJ/vQbY5L9B4U+MtX/Rt/je/RXZNKjaorMrqAOm4LDBHPJXZ+PPeovxsVnHkEJk5QqSAbALKcV
/a+CBm1IkWivCFycfJVpw+eRKBC9johpztGxDXbd1vSNtrnr8yEE205eMUaIwxmjwVm5+u5G6nFX
MMIfh+MmNaVRIpBWn7H8HeIfJ7vExGBKw1S/Cl9I6Z+9/tOxCV406tq2XZnja72Cq88YZ+nhCsrh
bxpjUbbIxBye7H4TUoP/K24jahN8la5YzgoLQNaoh3braCnloszTM/4glBr/+TQB5lUnutHW85Py
dSA0kX8sp293GYhxxQGzepKiUABjmNB/6gV/+83deRZbJlhxnpDDdr5LXF7dAhrrql56PtOvz32b
NVUYNXdYjWN89TxJjW+4+EyIbFC6kjDzXzufiwv71iPOzySioJlm9JC/aL3Pr0Tmho4CMbbhX1hA
ZhYCYXys8QL4nRf4MsqXTOYPFGRJS5rd/uuR2fxvetv4AHOqNgVb1GjXd7WLvdzm3Y9LUjDoKCSg
BrkQ9kBEtyTvpk8tB6AjZ0Wa4RQ90ZB5yAwz2K+4Pvno44BQGRHCEu5fnDjg+hzrUgD7KOsUTXvv
qM/MSAvFFDfV/wvOcYRlBsEsEl5FnXRRNBSjAg0GJRLL+86bJLC5ABozF2f/53xWLHFwzf2ARkp4
Zzx6btgYYdcWgUZGpbBFPpnsY7/kHVWimWvW9GBjbhv0hS76F+kK/bZ83l00oQ5iYZ/NdAumxw2e
n3StsUCvMAX1SIph9olG8B8LyogtMoT8p+ycN6Z/56xVbmlvovViozj+kCDgBRnq2YMWWanev6El
wNDg55ecdWWnJN9V8j22jDtKGohr6haHMQvB+raW24+LAxaj+5SURlCMM/kAGLf2dFOwYSQjRTCk
i5ku/5zpkT0bqKsWW175dp+Lih+0csqQtPbCnmL4lRJbEUfou8bC3nj77yo4iY7SOv/SOJF12gzM
hQGk3nbzE1nlpouqkaNRyQWYpA9+0aS+UgbKAJvmjVtmHwn4QhdDqdgrL4KPJOMhS3vTpoCa/PC0
7fZtPwuprmp1DlDtjbzoLAa7OVNrStNdbCcSgy8FOLjR1nqRZKaLBKigibkTwAKve1FOhQHPoqSs
zWraYDonY5oyogiwxay4BcqaX1X1l0BhCGkdZ7oXdtp7DpepLCfPGDED/hmUAt8zMxxTMGQhRxhK
HmXzFNT1wAZ3qhww9NN2XrnzY5ZQO2TkSeQ79XWQnkeesKyXhWuyeZ75H3m/2LiJ+VnpiWKl+Igv
gtzR3ZtPUzJI0KBcolxxxbdRi7z8mCAw4LtJ+vBHVkpcFMjFeG5TfADmyGaT/EL3GVCBONSiqv/q
vMfZRqj2ipbWWbi7gVUdF+yhzwZNEg1QlOnAXURpXJa9GYZCphJs8PKlLwD3amE8GtdFc/4I+vjb
rPYT2YVTCsAcLoqAaEWAYYS0jqmihJ9T34Z7NIU3oJftG9H1HRzV5IRxgaMeQreM35Hj5U15k7KY
aBw287wk20oT6TbN3XgTREaft9p/E2cms3La/0RUEQ9eLTtQNKj+wS5e2gUnImEZqKtkFcJyKVR6
W7tWLUOhj99fHOV75O1ZetcmW7j/lt+AmgFrxkp/kRHyr7rSju1VQwG6hSb4gVi5pqU31MN+yene
J7i38zKz+HAWew0uhv6jv0k8G74VtjS6REkYvJK7AvQv/b/FEhCuc6XULzMdgD1N78U4lEBHHuul
8bvEzFH2kAVR9qVNld8ndrcgaSdZe8Jgh+S3b5XEJu3+RBu66f/mAzidcZN24jye+2dFIi7PtWqA
9ZQiMLSClcrSXZ0P4jITuAzZo4hQyntckXlPvX6Wpg19PFNgRXRU3w5lDOUE1bYtvtTKg02/Tzxh
7AlGdk1vVWgMd8f2eW3mQUZ2ZrOLZf/70/oh+/puetUs/QYJb07d7RRLQSsEJwwXKYXoYDPMrWJs
7tcRf/kks3LxhFmuiK+Zibi/2rlNocGDrnxrrKym40cbAIEY8My8wRYJcGX6ZIcfysnV/nibqJRp
JFCi6LUJfHucMXW15q8GwlCJS03N4lcOqo8lmIs4oUTcSRcYJnboF8MdG0cIt0RqseLYtNhX4m60
ucKIxunn6SkaJFKKWEH2Wq6taO5EZIl1sUgPwPS3D7fK7RJAbtZre95PSW+jDZcDAr6QLOpBHjjc
x5J6S/YFWAfHYnse49YwWKE3jOMGik79L+uj9QmmD3dExJSg/ENDMAmQ5kJ1F/lmjTR/088JvN6Z
NUc4mE/8vJbMcy6zUM3sbZSxFRGyRlL2B7ls0/rWQmBmh2PzOsD84rCjXuaD/arsxAzfHGmi2UT5
DxDjmujyhVYlQz4WZ6pQo7bWw9TJ0jvI0oN8IZeTVDBfxK5f++udqQxtI8HdTrde2JT/M/g/r3Ox
SiIVN5mXo/Dcy72MvorjlAMiHGbKj03oPveh/41H0Cz6ljv95yg0B5YTDAMVEM+XZOyOKKehCRfJ
nrouJ5MdbzJQgdmEkedPk8sAZldNfU2MIsLxuGEbFiimAopuoXRZyctJTMSosd6wE7HpEfh71fb+
v8YJBzumhHn53UtHkNJjNdjcfB5pMaTxQAnc4L5I9cThCAEvayUo2fHJoPvaSnGrCfKaULHSfX81
qJjHkx3odflnPiwYNB6/Cy1HfCgX4nqv5zNY3cGxxRlgQn4sLxKykgyIr7khbOu7fTfXbqfDnat+
PJA0pQI5WFj/H7+hhJwNtVHI8PvICzY1DkqctyY4gpd214+JyE2oG0ZsewyISg4iSphvUrx8n3ME
iKAxsfPh5GJ8WvSQkaTsTbKyF86yznv1qTkAC8c9AZl8rN1v5KDeEALQRHWqWZSS5ei1r2x4mht+
iEc/X4Pupfj3GnO9tAFqy2X65dBsyX3CatJHie2F1Wgj/HTmUJhDpAvJBXnp3Nrg2HqgkvsY2AT9
RFem+LfdSMwGeXmmq7Mdx1kjcYLG4zYWLnIPYGlKBGJHK13fHS8OiswviEbZW5ITqDXcuKeoEHc2
ZXDxY/QGIBuxn9NOPpH1i18GDusQNIge672eAZ6fHH5aed66/kPj2HvkYbVBtymXxQjlZiEZJsqg
FeaeyYaphY+4YI+wu3iVIkSXZGFfE5m9aqbTgNKBCVojBFaZDdKtTi9zCvWh1ykuda7/HKjtKvBe
JIxfOSz4KtqkjzcE66cnvzXDxA0CxnrIWrs/vY9yRHMY+fzp/ZYReHCr9WV37pfkRV0zD1+FRf84
O5krVKOK6gtfuep/A1ZIfw4QiDphpIagr+zQfiJPLd7cEkfUXVZBzlqIFlOpyBvlfS6x9l+c1qws
BDtBGCg+M99eHYyR7u6Msdo59ykhhTWQkgT8QVuvMFRUijhDt5ctIBnt3zAOg1dE5//0psgNwVuh
GMFvit1DE4Sam1SbYC8C0Rfly90T5IctTYSEcG8SrrpIPFS1fXuanZhQrOy3y1bzlwIwn0lMMMmE
JHCsbjjnBuEYZQyDy+7m5GTWDF4jFP8agRoy33x99AzKm61Cu3xebvav2KNxELPAcsIZn6BeCAyO
gDDRlMmNQ9uBzaPhses249TMpp7a3ToW1QltPDmno+8AZLCDPPhFV9uPeNXzVLmKH0hVWPLViuia
g5zoW2LHzJMZZBzzcasONL2B+miRJOdCvAh/Cj4t4ibvAQyUuomG0iufJg+HWa2YVxZBagf5Uifn
7yGYcuQ+htoTNmh/paMkVIjecLJbbLaUe1/jdedFd7NUvLhyKonPO9dtGb6r3OtO68yXFSTLaaF2
xTibgOMDgd+buYWH0fSgXuI+gQmdlwKDEN2gowLb3BgqJIKuhIbCRX+jbopLsvvjR2N/h2z9Z4X9
ZAdsffRnIQQLoFAraKtFXyLWyd4N9Z/UhPJBYBmvfkcuH1aIKY9GL3z5bo4b1CRyHz8c4w5JpJMj
UA8hT/Kmpn5Kh6x7Dt3+DBvWeUGJwYPfwH6xuoaY4Lo5e8tLuUBM7XIT4kpHZ57tXt2rCmLb80Wz
+nC/+n86kcYbz1dPIEifMIRXOyKlsf89jydBxgdDSBFiDEJlwVk2vtik49oYMkcz+sZNFxCEWNxO
kDrQwqLeLCf03HKLXIC+WqQGSXDKn3tS8iyUHZ8Darz17pjt64we2LeuAnLjfCSRl+cdbkLzwS3c
gkciXh72KMwy3d8rTAJpq7FTjsTqlSyqIP0A3P3K3HZQ00Tp3D8Po04LiFv0MBayUIcIlCE+Ai8h
jpYr/PM22qp5nEUtSZ69jjumN2SAaxydEhDtZlIqZ3R3tmHKkFSDcQi/OdarMAb3Esz1mgKjFzZU
RQh2FNr0lR25Sgde6YdGofTdU7YRSE1mvXAizmgs41gxCysUk3AdDvF0M0SOXsqm+aMC3ybHqogE
/HzL7XyINjSh8BzCUtdbmBm0tApeYscSnZJ3Z+G7AOgbAHX20LDS8yFjEQDj0lh+SeOgWEbrZryN
Yq32peR3+/tTeqdiH4wXaq9/AZ3xDMWKMN2sStyL0rzKkdGLJPq4fCdyxwnWmG9zMvDCJUDLYTbL
cVPcNIjKV0gbabKoewp9hiiJEmKMGu8rLWHkcgkRZ6B0AotCOKhqKS8Gtg+xiBNoSdOWCQymE4m5
RPo+bUBAa3QwofY62cuFpA2vOLP/virgZlvt52Etn6t008TemzTYNMJ36kujg6xxs6pM9uY1ay4R
pIOju68/quWzu8SBR5X+Ahggf69JnFhL0qd2OXyQDIbdcyi6ey9PGmzMD9g/bFcpFcMSJT10bBUV
EkmZls3ZC9rrhCpDzNda03YoSD3748DM3FWHMRF4dFDXoSDyNiBgrsxkM95JjMSV2wgP7tK8VpO9
zkwmb6PnfFCauYCen5oI5C7FpexzSQ4f2UY3OJUXnW4BKt6yj/u1N77vzOo4Vygx9+kEMNkXZN++
9i7zk2Czufu9v5+Is9V5WmoSACbSsnJyBKcNaSXwsSe+OZqtfGqi12pKs0RdYqIuCHbw4Q/LCyqd
Voy5A7wtYpqcoQaGoKGmznlkwCvdjRgZx05oJmbVCDlD/r4JkDvyJnuEjqmkgIXgjeGJdxaTFbLM
0JlXN0kacTXXD1MtJp7Io9YlBHGTt29PU92Trf9O+vhsCr3jSIXqkB1dpyeU3KsVOYMcI/R0+P/N
2Nb5vTL9asi3fKQE87juvOYEK3DXl048yLgJgY3rJJFxd/bSOeFXKNm9zjHh3SmFUg6o9rqHsP/6
yZJRbJJaoNpoXUvzoPNJzYuH71PhHbjk4kzkOVgQq5ZN5KePqugFc+h2+TWT4lftqQ0tHj0yBR0M
rsooUrG/RyOLG/jfGmBRZG7l7PbGmvIRIBLHEKrXzO7HX6FRMgQBxEmhsT3rJRtaMSeZcW3Of9Az
AHaO3hr/1+lOae7FD9iCsN3si4L8ViRQvtOn/Z5sPYbSHe9YSPAIuLyIFPi1G0Trh58XpSk5JtYw
kxoi0Xhrf3czqTjyZIIgG66UrMLWq59iKjW6uL9fWBTcy8QTw5nV24DwbuAny00q8gE06Hf50q0R
8JDnkGxvA5gNEBrzu9Q6E/TxCtKXmD+kj6hT9QROWV7+u3EeveVz7P0oszd22w+bm1M3aa8Y+YSZ
UNP752cgUjQtUABWN6oy18rvUdLnKH/eApWrzXnZCsE+VEApBAGq01+sTIZiPiiTMKri7fD2Gvqo
zFR+qrlrJvqpSF6XHlSatkTvH0/JMdEO3Orqe84kv0uMJ98odeWvvg9jzVwXWCAzQ1pOKjAwcFjR
i2duJO3A//WzczPVScEnyRm1B5d/WqLh37S92HM/n+LaliAGqqc/laSw+HqCRA90zuakxRPtzPV/
uk5RF7yykbJrbn28CYUuO8ZLiunlABZ3Vr1YW5PH0N4L9FzwZAJGSvcfNGKWQyC/F+LdO4wzo5+c
DH/sLmZjk+prMmmX60x6aa0jI/EnSJoFYaGaO434gNfkMVlX5plYaHKwRmMDzCT7dr9T5o/2JM2q
Zt8cWpuEWD9zWPsS3JsyIri9wDUpjiR7tMjsk+4Tmj5r0OmJvvxRrY81V5ywuR375PW/rlLskhlx
jEMgZ5OZnr2X81gZrUnwy2KzeoZRUzm8yIdYOS2s3+jVPOBS8oMp0v5HYcJ7V7C7MLoZ4SvyHh3A
leIrzlO9xlWhSDX3/DKbo7n7d0oXgmvARL89wNJHUO4labYR0fiAFtv+9FLwLZvEH75DLqRSPLlg
xsCNB3OwjAv6LNDdc+rscWyxtxIquJrhRx4Rc549pbBg09XGOX4A98Y6nnF5IIqrV6QeR8nXED8N
fR3ybR9/1UQ2sVv8tcWezBV2T+lqRkFdTffg9v8f8THUWBDx/JnS2spgKi02t7WhRX1iSC/gr4J8
etyXdn7GBQ9h2DpB9oud9FYYlJ/q6khwo/+uzJp+jYTC4H5pbHNKI08Cl+nYBF09tRYksks6Hq6Z
E2F4kG5YGijtk6Cgno6uBpq6TJ3X7ZImOuUDEn/1DGAjHshDUNGjEb1Rk/PWX1IZ+O/hpBs5Crp+
MY6OxFCyiXrurBNc6G75CvydErRBbBrC2bH49GaXJSPPX8aeAbOLP79ukdSSWdgTqnj0cgG2+NbA
1peEXZ6NqH1mOIiluSwIPDN7lhAIv98Go8YM2edzNQ7EBNdYNpgPt02VZGUR8qFQXOB2PWdiQadx
8Cf/OCtFz2m6IzTsdfEDfJakD8LprDORO5baavwTWyvxuoLPJae4M5ldFCohp9vONx54NkH6nkv+
IgbQgDqA2F47mHzEoroM4IFuOGihGbFiOHR427w20DHtcucmEywiaQ+q3HIXqZy2EHPKe0KOl0iW
NHSdUf3DA168bF9UTs28evhNna2/PNWhTnn04FH1ukkYmKWnSOKOlH+wgA5y223i/bSsR3zEQ3lk
XqSWRsLXVKncBEh3dSFq4HFCUWRP8nuwGBgF77p69puM92fkJqoODD+Sl7oRE5HtNR7elK/wBB/i
mO7hy6i4lhsxt+wp/yiv2RZ1cP0SOfCu5IOlFpyaTftl7lPTk9DRKU8YeVLCuof8OWJqbVPOZ3HU
5bEQoVnrGG93BTC48h7a2SQ8BScCAyHiAQ7z+Qp9S3wGfmtL/tOq1D6VIEskpdBJiJGZ7PW8CbAO
hGv0JroITbK4oPgd0dCcXI3E60YlHPn4hvpV6PuYtR3AlWFFU0JzwU0/kOuj1KS7iIOINhYMCM6f
/VsmuyTuz/uv0u9uvU0Gz1x0yHFERK3TsVkmsSI9WTPNZXqOdFxxOnaQ3cy1xegKR/Aw4igoDLQU
DTuF9UezDVzXsNgEPkIZVYeMQ1dy/crqGctsVZj97/gi2NZ1VVuUlX0Ym+FVvruXy6xp7x6HEORC
hS//p6uroz3GC2qxLH7HqO7N8g3zcWb0erfJuvO966vpelPPgoQOuhJgHUAgkgrQ5VrRQX+EHf8R
zRGr3tZIyEkkodHcQ92pCr66tUYVXs8BXNDz9F3lY6v81RyK+GWQoHK8zLBoVvB4oixrDk/7u1DY
GpsxiEkQ7vf6wDbRfKMFv4doAjfbBBvHR/IcuG6GvE2w5QgZ2AMpCTBS4zcuFplBTh94fJ1/zcAT
rHOnFHc8NZfl8ApQnE5xHZRaPdZIRdQhZl96hx209GPvAERMhyMdFd+1STfI/A3pC7b+OewagMYC
wpDF8eYgAR2Ky/WOWv878xnxCSFy59J99yTgM3Zuvjq0p4vAMEcTsrvHHuxpCopWKoHvdjeMX2ls
5fhIwC7gusFw64BVZFRG/ANNFQ8ekClpnbUqIqvOx9rTrfCTYUUGyjreqrPVKUIXV5s0hDIVbASE
5KAOwR25ggyXR4mA7WhTYgNTBfbvZSHimSZQ3HNijLIWaNnoAK9oV/SsO2SlVre+eTX7zgp7FVfj
NMHZeBcwnB8vTI7AFFamrKpllnhU/UWxGUDe3kyzxKvkMb/jJ8IuiAjmPVxl3F33XCPDQHJRHvRk
AH0hE/FOqCiN58CrnyJ4xPsNsA3qgr5E5zShmSG00Xf8zNYX0xM+535g32ZIUEUK/inQkNchiusW
R5acn3sJoXadKc9n5XWiBRwpnGIpE80gXjdGr2XRG2uBKc/D+wGpbVUwUhV3iV5+/7XpC1t6sb3j
cgpiedWeq3SjmgEtzD7eP/qr57vaBo0pcs9S68aqpGZw4t97AvUnHsLfGpxxHfDfVExYqN9hu5Vv
IclVx5vos5xgrjVhYPq0wivsp3X1q+6dOhsQHhni2CPTr1AICzoEN4eVTH9aSfIGdKOjsXLJ3cJs
qFVey0vRQcTyEV+mNs2LupMcAbuI5uPgDsQHqiHkMp8VXkdFhRaSTfxyuTym/d7HdZRFB/mQPeD1
aXmCzLt4ohqQh5OVmW6B29GHLqgLsunKTQetgla+98dePZ85fHwgjQkGyRi0iLrc2/op4T4Ck+D9
/9QSAoTbAw1PkPYRkGZCchwYwAlLwbmD5N9egeMYImKx00z/su7Hm0aVEJZ0F1em1h9lx3KqroH+
67BBJrkWzRSXcBYnEvLeK8CrhRR+Sllytww2zhEThf86pdF6U+mYSPv8E+m1B7paDa5CLOLMbfe3
zaSRBIUnEvZyoJqt1RUzORJc0PZ6Y7mw/dgC8uiNexCrAHZ25R+3HflGEDwI7BMnjpuGZzWPlDpt
LCDPkZL9eX1wqWoL/R0ZN2aZKQQhQvrJM4hsu9bSup74s9mW5AKVL0+AeVPSq5mD+QSi6P5SXBsB
NzxPaLvZEpWIUY/B3Y5CGuAt5PxO6JpHTHfGE8Z/j8gd2nXiJ44I+xO6PGFBEcbnJ60BgP0/43Nh
IaDh892b3/vqhKxDwZ6t+O7XIOQH7/zwLGbanlFXWv4+TDqo0kcO/HEr9uo7DTYSfsze1XdvRzG4
haNk/+y98ixHaiKInE8D0xn+npN6/V7YZkptCfRfMjckbb1zotlFdy54h/2kxOYVCRCYwjhkkWlZ
JxeACleC4Zrp5vOKj0OCtER7Xw6iHDV1DjDrhsPyVnWhWx6jf4s4dYUChNQk8TEhNofgdJMt1unB
SOvZgrFQJZsV1U6DcoF9C36QtmWXtTCP+myeFaaNFpHkaPakzQFXXseqMj/hKfIZbIZZGSXasHJA
9Ale0Z5dWSn236KbChPmP1Yk4ONBPv9PfwlWmJUElHi8iN643nLaBbuk495nczUegh9JwtUdPqwL
12zoYLu3tDtIpOXPeGkcJvc6AJW0ZtXLnmgLPiGEGLDTvLDiedBpWyVPnsWR+RQE7NV/9mqU7RVr
4aBKB4jTelX6Mn8vbapjkbJuM1tm7kX0oNiP+Qme+Uap/8VI1MXcKcUbHMcmxz6CY6ZAYqViBGTe
WEFvGGdlvhQyib/8dQIkSBN7EQ58BcFpvntDQqojcSUSjUiboljsruhnSuZS4i5LOD05FT68uz1i
aVboN3n60SYPCTG+kSYvmyb9s6ROWPo5ApCtcnbds/CIaMpAEZgNL6UkP3yg4jNid8rbtg3zCax2
2t/AFhvaqQMB5wSraN3b0Fde40d/JUPpx+xK3uXSbJN24B8/pdOCD/KLU1kT8KI6E2V/Dbt5CZPB
k+XCkSM/UYkAqBVeS3ed+yL99nA90ZWzga++VQmX1UP0u+tNg2lNE78atD4QNc4ZEo5FUaaOI35t
M4r0UBit2EsudMGdEwTp0t0WkI0hpl2k/9BTp4srmFYjXNlHnXZ76dXdseNEyTWhZxz/R1AQGb0s
bEOlJArXp7en+v+BG48lekNg5lT/xUmI5/qQodF2AOc4HqVAyEzb2QRO9iw6ugn5K+wBWNefSpWq
B2b18hYpPfV2g1AXxJ6O/P7484O265nd65yMXc4Ornp9+yadUXYlTNO4PtVNBX2G6TeU3FA/F9Q8
iDbmhn9UV1TcMHGkU+zPWMbutZmXsHbcaupUv22xlXSeJ9kUwG4SSdkIJuQkH0GlGN1fiLY1TLSH
TmaKXiZJAB6Xo2+NZiHl9FDfhwHj7PiiFyzT2VnNRa0AkxlxQ9tX2tn407ItmyJTEuCZWw12sVh6
envAwaF7rh6qJQgM8G59u48CfinahJG0Oact7YmmiQrEh9lRIAzK5zfyFbAjuIpwBOuWgxcFUh+C
6sct+qLj/gQRQGyIwGQOAOFJ5gBxkDh9MBQ182XLO9vN/093rflrLCJrX4NqABypuTD8IzPtfxWB
QOz62wnct0ROd6OsV4EoSwsRBiMMDOXJy/4uAvPGCHCtJZC6gwTnkwIouH3iEslA5xqqR3F3sBoB
8ece4oi0boYScGL2kUahw2Mvk24PTCnrLMdR3uTxM4utXnH6g8SGP1B5YKTHurK+/f83MwTkjUvy
mszofWdVvL71Tl1A42waAMo0atJIZR8qICZvD2FYxlhWrw/lspj435R9Uz6ZSRiMEIRGfBks1pxc
rz8hCg4l2W48I7OyPk3vC4nRFHROUkOwIjJUViSVfOHhShaZgCgmN+86MDv+YbGKd99XeDBrDmuK
4f5K1Ivn6qdGiVrvlzuzHwNC9D3JS3pDOPf3/ymFhM39OrpT8y043cSlqCvhgSx2zTUzQF0VsDni
L4kdJYE6tSIUBr9BkOdIs2E+y6Qs5SZHDuv4NXDsQA0pwIidN4s54S+wDibiJCC0SflFI4VlOwB3
j7/WH+YHDfYDthqqBKCSyQjPR6G0H66SONlk1K4wi49FO8kRsefnxvX8QP9Rmn2HuOp4i8Dc3mC6
pzYNTvxIPcIEpq+TnsmIxJzDhpqxip4oxv6//GLiq7ljznd2uoCQVKRPLKjqn2+POtVYnAoKfKUp
vOU3+Su1lFzSbaHmK/lAfhJJkaPrhETSG7IZ7rvo3Gnn83Fhb7BBkBcdhSSrfa2JTRwd2CemBx4Z
PksNRyRoqujeHcRqOZSM1+hJrs89B7zl9YQtw6lAKpyQUHM7sbs3ava8RQPHiSbgcSN0me4jX1nI
HLFgNwVhHRUT+zgGZr8vVm+TCZY0n95DlLd5BCV06hJegFCxVji/U0REy/mI1qX2dmqEPHzyY5k5
YvBMCecrQhnJFI9sEOOkDjNZddQIiTpBT/gIY1WtZMyB6ha2voWvzSdttn6wNtZsUnwOlCiBfEG4
yBfEnwVwtvexWrQy6SyL9Zci1ARlxuxpY21us63f7dMMv1xbgH/AwR8O9xmILm+YlDRQ6Lj4EjsQ
vSRZ2CWPWX8uLqicHxD0crF/pyEHGY6unRYAuhz3GQ0CzkehlOzqyhSA1jV4lJFoV+n2YLk5scKq
xZ9dIbE/SB0C/y4eqtpmKOisPGZ3ivKcJWxtaSuowAyTHTEB5srPL5aFUk5NX2sJkgQDzax50r/U
gS+o9HLxEED69NJdfXLNUTqqRmbhh60//PQxfIPIKxTlJTUAmd4OVEd726NBCbuA3NahYIuTqR9E
RfeR9bq0bd1uaVrVGQI8l75t8Iba6zZLcLCKOHWjEsLbDXrMmwY2zUQUtX8PsyQfBvjjXwJomc9N
Y8OHIH3UV3kr2pJoftcNbEEciN3t3L3HSoOQPjcU2bHzgUW7co4rCuLpXvkIqko4rdG1X9oEJ0yC
G9JtsyhrL4TiAYV8cD0NQyR9xYab137sYH673VDKVLH4OmBgOsmaf4X/M19J5LAnrqs0u0fwPp+A
8TNTjyvoV19+xn9lI0/jr9Bx84VEgd+XsYfaKvtUBA+LwMmT4x6TBycSUA9PZ2Wc7OOvVjCiEo62
/mM9j8qfZBUJCLsy4vhKGVPkM8F+QU2kAvwLuFmfS7U3N0Wu18JPP1UN3DdjRNyXt7MGjxti/u0l
hfinkR/dfFk3s+ofsUsZ527rxaDy6Zw6MwElII8TmdtUTpulaJHaUH/MSU2ePKbER3Y6MMZOQ1GY
fAXoRToivpCw7rH/OipSgIt7txplelz62RBAnco7irzVfPnkY2GsKXSpUUODZ3mrK6ywFNx68bE7
HOE2jnYGYL13URAOvD3U+wKHX/2cdbygtMvlxDF0ROHPbIi0uXyZnjaZjR2rKdRUSNYn6RsPFEvi
qx7GXH4gLwHDO5hOBDnau/Y1qdFSi5U/V+dcT2wsnKYnIsd83CXiHJXPXrFv+usbuNhbruQBM8Fp
Ps6E5XoRwjyODbnqEWvZG7Typtiw6d4iOYJcv91P+cF4DXclds5fUH/6flDODtXHSBSn3n9K5VSU
df9EJdDYw9kWeOvg+OLMNr1pjpGWBORhelAuTri1JSIwipm27/EOBspHn+HeRMKK76+JbxIUxr2P
5hqVcQTbO05+w394uALUpXPvOezVOO79tAmFK9lPOVix3tuqr+JwYSMY5FUCC29xQG6yW6HYFH8b
AayKEGXFOkGKdeIUVQ8U1KkBHpwGMOuywi2Zn3QN82f9k9Z3m1UxwH7Y9Cg/gW/OtneiNtAbUEHe
0w3WJFdCpQtabLNILdyabi1svnFqdHyKBD8QdEuy6MTN0hTOGhyBXQluVQrLzay+hhrGZ/EZ85dP
N6S+oR3fR9Hpf//Scb1oaCC5PuV2VOZmO9iuz1jGOxe/aUhJej/svqrpGMaEvqXfPuu//b8ePwGf
cx961+QrmD2Fi8DrhDWBzdcczEM/LGu1aAN21BkebSnZNDNMa/3lyPN47fJwrEIUuuMjdzo9im+o
YX/xzIV7deldRPp8mxtUmUKOIhNmSE0gkH8NboBHAHA+VP0Abhv+ziTcPt7NOmCZZNCVJTuwR1dA
qNDBd0QG0amlDRwOYQqKXPL9CPx7ghOpefUpgbl2kLELsgEW39KMeFacMM3/cGwRZzijadN1xrmk
Qz5ReSOxig32M2lqljeLI/BQKIajr+PIeyq+NCuAswIMqtFUMZq/EqhEN5qBmywZqk1BxWLFqpyh
IIQuIx7eMXIHdoEeMvDEOExG8x+l4J4kVJqSkFwQ3GwT4xQZ/kbs+z29+5tBrchu8hadWWdMifWc
qbV8YrAwoeZPmxrmVTTBRRMX6X3Dttadt9k+ctHiFvExc2/hNJP3KX3Itjdn8nLJv/CKgCIJueDD
OeuQz+hvlfmtTvbdyUwKsnqUMQHHMWH1827qWzpnUcru5kCGTZzRRvlMugJpUt8lZZmQLNXc28CV
0ec+pri/8z858xpXHzbb/n4thDMOOnmELFTBVNKKaqGri5JFvnasLD2n7r0DTFAAvBpJDohezGcr
Jg1D15+/DwF5LTk/uklhntuoDx8qV5GMIEjuAHF1uUmoM/jsEDI2P4V5ApRV0oV3dsuqWNGtjN0Y
V0pRFFD9fa1oD71pdzY2VxdWYMFGIvrkUGAfZn6ajGJ8PQOismeqQS3vjuLhTva38r+0WghR8Y33
QmwdqpEdkCEjlhzG8OH0ztNDdmJhMjB6zBlrmUO8ViTLJeCSUd3o59Z0jw1Rvv9NnFCDsA9CywFi
9GcmWuzVfTU+PJX6TxYC8T4B/VInMOrj5KFwhhSyjDeTnihihcXw4GM3JI+9WkWL1eFndXnSBw4O
wf0kFTXWFJwO9hEzEs2UgIlZYjlzMrTNWMdG2YhKzqikldrSE2jQlcUr2SxJM0kK9uVayaZK7msz
HpALycb3Ux86NLYYf4H/oMlwt1fbnVzXjszm6IfEwNuUscwji+b1nWt44CD5v8S26Ii69NI//k9a
Rz5ogxJmqEqL78INbAwajA0YZCT81QdoQJP7Nq+OtOuyXVj99eQ/TX+Yzm6IKXOWbcw896/1iu8E
eCIi7fjqX/vZWYPAFqKtPd/L8nQaXQKtgaf+7TEAYWY+D9QKID0TDjBghgLJZLG+6+CJDrow9rR9
30RZsPYBLrth4/Z3My8+2dRptPD1k4VRDmkBXpZxJ7k4PUKgyGbeN0UO6PXneFGmjgz/RGrBVzVF
rtIKHkiWcQf7iJtcU9C/cL0obwuTHhVspugn36RV5nR4hMl5rFrDtwXm6lJ7aCClkfMd3SboRN/k
XBegrsG+wylx0Jooyu4HAhnzXsySJ32Jgm6SRsOlwnTGTjpYI1HD2ojqPDXan2xUTfVRHciRS03/
05T5Lox7igKL5Hid3KERRROvGyYqce4oLNDRUb9wKp0FDASm7u0zqV7zd5V3xWdfx+920YnRDcHE
5sYic8exZAcWQEa2s5hfLd+hyEdCvZWABoZZjavpRKAJpSdSOS3vsi9rZez0HO561QwdpyrKyVuz
vnHPPI82/48Q41xFv7I4mJbqUE+TuaDmEVQ5BVM9XlOBgtLz7KtCYn7DGx2q2sk9negFzNx1xMTM
3gJ/QdilmpQW2Z4IV8mPONcZuPYzAh4PB4jhtMtl8N3w6UfAbB3eyB417IzuZlHioundn610MO7T
0DwCc6v70HT+H4ZaUhJaaAyKX1HdajRnPVj9IwIzjWdHcUHg/eUKij/yDSfyNuMOv/Zh70zRoYKQ
dQiiVsF0nTSLN59s9rWEu3uTzIVXzYAUZR2mUsHx7+QbmJDT50kvFJX8U43WM0NLkMKxiIfYp+iE
4IEleYXXbfO4HptiUNEQOJwbeTkjZdCgdcgUHGZ1v3sjcmsKzIUzwYqmix1JgCIdodt3sEGEliLx
Wjfx1GELaAN05W00pinOKQrEoPXCKm8CDobhf4CLaa3CPTLDEIZcopLE0qW9/TPFc3zM/dkgiaEW
TFkLLvRUh+pIUVU0bITFGMti6yVwwXv05PUxhC/iFj0dcMcWCurs+wKWyii7y6RiLUeM0jPhF1gP
UIGYnapI9wPXGJ7JdhTAYXTeqe2Uksfr+e7Vnxgxz0Pq6i/ZtziU2uf45rfLcZrL3DTRl/By7Rwx
W9lAZu5teITHfqRFhbbCfuqX8CRm9GspCqHHWAnSPNBhhzn7Yf1+Cz6NG5OX7Q0o+ikE14svVLHC
mWOLVSTz6bv4cynzxld461Ok4wMtzEm3VO6+JwwPR8MxiyOmMZ6lYf+1eHsqLXzVEmkHhLIPDA9/
+l2IQPUmb8hxrxe4aCDvwUlIsH9cOr39uVcUUDHZuc9IUUZ/F5X2Da94yOxxfL5mCE1GMDkeMIkI
qfAPD4wOSlD8UAW2oMEStAor4L8KiIaw0xnYoCQeRUQVk3ISuW9TGEAwdvNsjTT9MCZ8bLhdOgD4
BnytT7CfRNBP97AJ+EJlUDnI5ncv1cJXeZ5+LR1dtUu1kTSo31ZY7ZlCbhTVdWehp2/rOh7BSoHs
ubDbM8tboHoHP4Ccb/ntjVr0IqfSK88xJM+1P28rJ+11bEYRwS0TN193iAPxeQO1VD7bFXtRzjS2
IxNCOUcbjeCzNupQSsm0Nk2CTqfGJ6d/WKh6oezomLVhIGpdcWExHMc0ONjQhiT2IYLQ1bx8vZRV
VKp7c85ouXGYtpsFR3EqobWz9gpJMzYnnh5xiarStMq1wExptnh6WlM2IAkAIZFh5JBUsA83HZki
zwiaJ7MyiOpdF9zF6pea3PUHlxwGNkiPzhj7/QoAxMszTh8c2R5rAe+t9oM9zr7WcoGx8ujy4RxK
UoPDl3PbeQo8GnuY67j0NgCU3HQBLh/8aIbmLM4dCOQtM6xz4XkoNMXC9+Jae51wszyljNtOirVb
pnBF52+KU2L4dTYgn97D/u8IQrBad61Iyt4HTXf88TFSIvqpl/7hsPIyTPLzXwaH7euwjNohgG03
S5/4fT+UCWdeGFzd7FAEOR3h+tqiyAGGG7aN2BSn7Dtv9/p6ZeSxLgkScYU0pqdzRW9scJyQVrcR
0KbeEt1xj2IWLNpcdluCsusMifCyueeSM7ll9vzNwf+LQu51WkHfeLxbtdTnixBZbQ2Lxug/WNDJ
HYxsslxr0ndN+UVeb7kgtFDpWjnb8sRbL0BqIHvEFxzHwKtl40wHjBmlyJBA2YUuKrZvTOt1avq6
vDMvYm1mQumRBvG/cAayKnH1Op5Zfe4WaDjx7XuR9flgZSS8JCwsS71hvVWH5NkR7ZnnZi/Vj2St
BvB2zs6vXoM4oRtpJsxUekKCc3jsI4NYmikPDAMa1tLR+0OtmHWuW/7YXRIPoL5nq1kvyYWDw+yl
PdtatpNd6CP28VJ7BpTpdOoXo8ZT/HyFRamZ/I6r0R04ATSt0N6d2L96jLaBJ99zd3ZHHSEZhnOF
iHJz7bJzO5fDrBIW7q3Ng7NLbTI9khsAsQqAIWy9O+eAqgEUAtJ56FpUcyWSMSH1R0Qs/UZL72wu
bd9awaz5DLWjRfSCezzqJ3+4YO9MNkXEJq+rdM7eCc8jjNHZ/0MU8bkF61SBr6etKyPI8aAgfjrC
0AZp7NfOJLSf6BwMHO3ckwBQewAzeYx5Yp0Vg2oq7mg1a8UlWD+jRdG7R3C+2pM8qDkDlnWSj1vV
/BVFMLX9XQv/DRQmwCmDvl46AApnAMopBIKo/zXy0g/5ANtDJumPops0xVbI7vUlSsxcAxNhR6zt
J9zPx3FtYlZSVDao+Z+B+SITXk1QQ1QCyqYZfaDutC2OMYIPkkE1XlNhJAP2yy8R55rSHOBoA7xf
rGeoaEHTkPZoPMjaRtqiFbft0su/sBtr1a378oBfA0zlOZos40t0QnS2IUroE7/Hk6PpD1fOHotM
T3xi6RkkXzUSsQJyCe5KmAjnDi4H0hHv2DEWJLxHnu0s/prNKO8YsZmC2RMrDZaCMMgQ+ZQXMD1R
i3uCegnEoSGC5mjS8P6c/TRKZgfjOECsferyQnDq27OHc1VUQTpIO4FsXseWL8Necy9s/lQtaGGs
6BYDcDAi1Vw+crX90yDQqKfGA4rdID1Wheg48030LP23u31+Py+Xab5RcP8BVWOs5T+gNU2ryN18
EMggbLPghQi6v5FjKFwwAdb8a9S8yhob886ROnpHMTslm33Z26czS2y2rg3ZTn0m1mUDPgSpacZG
Tu7grqNiF0IlfDh6Vsj7Ttit6RiNW976MrFi2ohrrgULD2bo2DfrAlTN9fmPNl1ukcvTIl3/+ocL
hSG0UnXM7SMbJJ54ksOL8gHMgPN3ngaqhfTOID8d/FfwwxuVThVfZn3FOmT6OI7s79FIoYqcbs3a
ELeRkC3O4p+zsOikzlGSwMi2L4XXcQNt7aLJhFg1KJBQjWvnhww+GwOdLtH/mLS1ss/q7YPv9phZ
cvLJJvbcMtm5AK170kZcAjFsT/TgmR/0LHnhmBlrHd7Py+LoYCDSzsmfI5+WdvAVykZuBk7Icpj5
2Z5y8zDgTTrsXqTCgIctLa1QnU3/R263+np2PHtwni6MIn0WSfr6iqQ1ee1xLb9La+YE71RADOF1
C4JPbYlFsariW8yp8dtNR7N7M1asMYSArvX3JruhPhyaAl87JXQBFzeepi/bleGl7IcCghGFXIMG
Lu1eg0zqh92iCMCAed29bDaWPxGVFCeKHYyDa3xn0pKZkWP/c4WS7hoYC3/wvSgmeYsnMWe18Xog
h3IF8HJlT06Ya6awbSQqkfZODx+lge37OvsJpBbGLCRXFWugRRvx7uOgfnPdT4R7vNY28CX5ZHSF
iZbjWYXKzE8uJsqolC3yfaKFe1ATE9jq8lQule8MQ4HtT5eLJZjogmHTpi4UewHzI+A8hfS564US
nVpFVsv3fFD4LMQXz+EDGSXNpQO4pyzX8oX/WaPjwqkRGZC9Ap89ugjcxaja27DjukLqmXoAooUA
XdtsA7x4iPRB3+aFNuJENBrlV3C8I++9IFT1cCUF5oiC2rG/53miihAG1yeIiCmSJEMnWauYEzPE
nPRnS0LeZAHjcowMMTVMK2eaJ08ACghaEVTpEfe48K0qv/mdW7VjL7Yi83fg1o0T2T9Dxoqvv0Jw
dY9Ntj6q5AO8S5D7G4+WrvdE/0MptEApsqJDZX0AEZBOoSYYRIP/rIorVzmWlGoixp3lQPNUb/4Q
LebMl/A+ORNud1vEans3yAdGyUDciB/k8oArw/4eUVfleN0s1InXAaQPdE/z6oV1sEm0cGh1Bpza
rR+GW2SNrk5BO9oBtAoXm7+OajM1xhkBngEUy4hMLUpH37Vjgy6dtAplk0Fm5dSM94QFoKZGlbJM
yhuUo6yDhlGuhqPnZ2IvslyPN2mV55URo6kCtGMb7szbDH8ifxlAPS4tLurAHIGyfoP/iMkxHlkD
q1IRx9Atj7CJ1HCxU6+92LRCCyAGj5oQKP5iAT8RYI+/GqwBSibQrpwVIY6fmWoUJwy4TTSJiIVh
sg1fJZcl/zIuGi/2rreykItBWHJEUrs33B+NaDdOYbug1hZEWYou/8h32Numd09ku3PqreI+4SRp
4Ub+L7hLh36x95+7lBcC7gCMl7D2xX2n9QN9WZbKm4HAjatNWxHp9TxV3xE1PBQPm6MuBtyHF8td
RY8Tv9sgXinAlLxOpBe6/6lL0FvRgBBWUF0tQVc8Pvm39vNSK3GJp4goCyuw4joMmJpJp77X6t6X
/rZ94qjiQOZlc656IPCnyDO++3RkZWCCAZM7xq3Z/7C2MF1xand3DEehiq8wA4tkCf7TfMhhJt+1
kHyfIt2pXmZsCpaMnB8Ef+cUK9qHwe51lAsiuSEHw8OZmE9Lv/s/fyFTKoYBAVryaNkKf4ClJNrm
7F/+En9NipbawExKmKLZ0lfvfslbKM/guHNCOLWtGU1bY6A2KRSg6OHW9JAwIsmL7xBDemzxSGry
uBxJYg0oSa7Ho5DSNTotd1L8p5m8oi57JJlBP/ADyYjsXXnjIxS1MVoZOBcsflUxhBRT5fR2k5T/
a2wXVxYGEVT3UUZ1qbuzUk4xQW6nnuRdgCBktrWDTrCfVQ3pmgxJV2N8bquV911p1abL86t3eJ3a
CKumQ7jFuvT4K4+f6IUB5gOUoBwgfU9G8DQywlUFGqG9pOg3YYS+e7ZvveF9gUzpcOUxZvadTwAX
Y7Q8U5PCIRMqz5j6gdM9b8GUUe2HL9u0+ciIj/mlmJt0MoEHeMsWR4QszCJAOaaMUANbhiyfbImf
/4QXoREvUHmkmVX4VbbiL8j9EwG2nYOpCgvPgoa+xwV6MEcaZebk9remUPbEeyjM3ZFRQHItIC0t
IqEXaav4fLvSP1o+hJ+hOtpEwoMteVXWV+BEVUsIUilgmYjldcTAkkz8Tc8HMM/CbNuX/CzzExVj
psXwfFbXS5JiwWHU85DdoVtXRW27XSYFnXUOGEifXdshEKaCR/GJ7jWNwoe9yy1lyHkr9svl2lsa
ca4f9rIG+iq9Zexmxp7dQJgI851KAGiVmP28ngB2beXZpa4+glSxM50cJGXZU0nFFVBxGV94clXY
9l4oObGryefW2jdYxrI0Mw55scmFIkdWixPaoZ5koCsrhJwcme+Zc9Lh9LOBJ8Taw2FkAxlPy7Ml
z95i1+1CQtXTgNfcvvVRgrrT7Oh5tPnPWFGIEuYAc6uz6fCMvnkk6wfDWrAg7RNnoajIFxMXnHKS
C53ec/rqEhOZHjIFai73CibZkH+hBoAOFY1zda4UT3yMSSwKB5dQxQzOLLygoPV7weCs07GSTFox
Y69mxcD2a1CJV3j/rT7dD6TUL9Y2/fbhDqwMaS7ytI+d5y7UiYY3TpFEtygaK2v72/xXwjDGKI+v
p9/oRVmMSsQ4jDmP6VGogziCUGtaTuaepPnP4++UJI8XRuuJ75aiqaX4cFwAuOvdY+O6eaVcYdR4
nl7rh9MJc8v37RB9D8WtxQf6220X4/d68XaKu+wC+U6jGBo2R+zRUG9k3yqjHXUWk+G9SQVw3+pp
GoTn4SQBlRL9DnnWz3ZFPAPmlpSXWp1N4UHa2j/66b8jEH70wlMO7vL6YXKtpYO+Eqk1rU16kqnd
rVw7oi5XRKLGGPjCW2VgLwu+6bWrzxM+gyixyYROsZ2f876Mw8WuUSweiG7zk5Bu6z1PDFQIIzWW
hJg2TDVw266q64DXgi8dhccY783w98LeyAdvmovNhgIRY/vTkKoJ5oT57tdktWTTpebXSUWPI1so
1dXeM/Vr6qDoCnaslJUBn8rF5vao4Cmj9zpd+y8DE+c5gKRB625TBMdCONthkHW7Va7hXUA6y2N+
Dib04JVtSQP3itrURh0SRyhojCLBk0EnSkWpFqLWXy0Vmlu7PT51qp2mfVvaXqnManDTuu2UWRGS
O6C/bgWGYZmGxNzpH4cyD+gK9Hs2DIPQxX3gRVAtbj4Zf1VmvJNBg5yO0ycfXtuDDg65Ejwd84qk
RYXthlWoIQPv0XXI3pLId3Lta6KZ04TmdocMQ/eZeYeNtBZyyLjSxQxWjxtkfhaVCDiiFWVzyn3+
ccDzpnbUwkWOqeX4k8ZaonleZa9+d8qToD6RLUVbssH1KSfk+bu45ns/P4opNpH/fO6OfS0x5RRI
3rAN56Fx/JqmviWf4vdMG2EYb5qRDtKrM+HpbctHdswEaZgWCpbFnQGzzTpn+dIi6yNlq2THK7CK
xyHvPAQrE3NKEtN63fCvWq0ir/NuHmy/Iy4zeCm/H9a7VIcZRmT0RYHZKhUEsb8mQGVgQAQ81+O2
WdsVJf8mDnU+xuNbQ5UbvvOu73eYwnpAXo1qFEGMw+On8v6uH02uEC4LU3cOcFR12x4gRXVE671s
i0F8N9umzLnWC4QuooO2KAU21kdiLenBYfkxpSJrtoKHhGC/9XqQus8GkNsPrIkZI4fwjjoMI0YE
iBFdxgOjPWgUi1zAkcp14tzo/k4s7hzWHTXNB4ZaBCcG+oeBJFcMjjCuic9ReFXXVffO3OYKvpXD
xPWiyNH/l+gPkkL4KVC3R3VncgnRLHSa9olSk2RWsUzG+wdD6NBHKkBI7osyuUz6lRGpo9kumA4I
8rDJkT8LoyZsK1kHtd2M+1ZgdlYQBg8x/UCCNnDRAHUDANqfqQT3Y7Jx2nUcroW6OzZ7VDQNmXDM
8Zk4wDGpQEpnZ1hniPbXxToDjbuAHFjT6VNwu+vslbFRvZ7sWzGGjpNGtH6ILVxkmuzsIFKSN+jd
vnl/RT72ADB2+OVxV/dESdXzwr05Ryqc8szL4Cte1rLaVJ/HDrFW+aVnk9Yv/790BfLPhXBNn75b
I4TzAMVw/DRH96JssjM7c5Cr2ImQ9Uf9yrDK13mDKQmEybO8WZF0zGusLoz3whkePTMoQ9WxGYwT
iLbVLjSvFI0/P2uVLge61LFhTNpeZ7QeZBQ3qf8Qlyfr5neE+CfKE79t+0p/RWw4XGiHebAPlV71
DJ073vYuozPC0yqsp0EBWlW0HcnSkCSNtcgGYYQNMWq4YP0EBlIU4ErAPZWwUjb9F8+k8SI5wnCc
os5h0QgMQQgJ1qLWcI09OZkoME7YSeLZHidguogYvpPcAemJYeVQeB5BS3Q75bNQNNaE0YH2X0QG
LZWUe3MHZ8cisj73geOqVOiWfwYtGKoLZtIMagrqx7u6Db94Tz4wq8nZZysS5kUcKKrE3Lq5qiAh
hz//B8I66kHpBoXrNCJxGgtFeI6dfG9m1uD//QCp38KgTsF6i//UXxPmpBIS1k4XPjihavgeSQ2e
XKaWbdEJP0/ujENgFG0uKeib7uPw3zeXG8czgUWbTQXzVvikKnf3IApAwijpWyh1gledwdXGBfgP
m1Msc/U68ELwZL+iG0kTTbYr32dGOt5xcH6FcGVmB3qujwg0XMc/WnTT85f1dnMAj1BFXbLDjw1Y
QT6O1KbotGnCQK8PYnHdNqQtwTZG1kl3RHP45VKEdyIVjK8w11haMFOhnzHGpz1cZ2Ps9wKc7EUj
EClIaVzGZuAcYWn+GSrG4jB91CeKe4ycNRmQetSiBG2ZpID1CmK3279rvgLcMzKHVi27+zh6aRjn
wSu/fleoCeDfcU0CN3NOToSMwtqRwQ6c5gVPH+qIOuJB98lGNddfpCesOSSJ5uRhOU6NS7k5PX4I
aVwnoKtWob1rkDwKC1Wr3wcifIXzJlZUyIKQ+IXYK0B4CNaZV7EDfwlQacXQ30/3/SJ9ABEfieis
gPtp11kkRh0H4/8q595V8WUXFzk+vKuEf1+d7393cOwIna9tCgCL/thPiAz1WCoQ6Mn9SZD3z1ip
Q/QggcxA9/jm7k1NKaBPCdfJ7itVCRYVL6T3Tl+8KRRpAPM70p3tKaJRmuf/SYvDfpT1thWL91zR
R2KDqWY0WcztG8klsC6Y9SLtV5I7bvR7uAo9japqJKAr9S3n0CNP3mCki0anWvtVblR3l0RumJUy
JDsrmwgxZBcQVGI6ht7QvV7LQDI3A94/t9D2VNYQqOxXwkHu74AwL2O4vR70XUUfQkJ18+s2ug8I
YJoShZolaT4dNKfk7Ik1XnHS+aaD4Kkwp6jLlPmCqppS+xADlCUEj6J1Ey/VJPiwpUDz0VDIM02J
Fl4y4HifsoVfuOjojs1p+rZKi9PqXSd9XxHjAV0nThwUq+vinYZu9vFd1bxxdN0nDutxBt1TneET
eweM80dToCY+tPNPpM30AQw34LtUTNoXj8H8VeQXVhYWDKvG2pwYAtW9H5Aj4ICCL7eYyt1ZJ1cI
d8gvjKkbjTwtjOZijZS6pRLMug3rrKn23tSLTslzuDIhSofPuQ2GLuqOmPkPB9fUcODE6AEUfOAG
sSuoCPviq5/wOlLFHecV3FG6QnVOeHzS9kJTX5aB71rEYtS7acK27ocu+nHHZ04808zMLYuKrg9T
n/037lA3Upnb8Qo9NXEL+Wv9egIc+DyMi0wM2IRBs4xn8mr6UAsal888rSW1Vguhy5Etqra8NDmg
sHppdOWpIr1ufFBxceqoX7VUoem4oI4KkHgie4Vu7qz6fDk70h/Tm0mEDaqtg9UvTuoV6qiMfV34
WOPEDM+kowoK3/nYxLMCl+KJxkKNV14qeNLg4lLux664jG/fuQL3PZ4wR/K5AhmqpMvo2BqOHjCm
Qpc/QmZzlglb3r652FIvEUvIQ2gcgl7YHs44ooZXBo/bhKno0obx+Hq8/jDaLgz5AtwklrQygFKk
BLOCq0/16x7HU3CsQjtuQPsZ3uRgJAncxniL52XYdpc4mLALJMCM863y0UFrV32ZZaAfEYtmdsw4
+mXWrmL0LQgVRGJcKByAfXdFnP57FxMe413sbWY9+4KzOSMLIGNs5PSl3iREdjS5U2nxjSG7uRy5
H4ih3qBVlmPDcpGXB4MaU6meE8bG/bzPSIrQUupyKUc8u5lgLUsCYOIZ2xt0QD8qX8KL6vgMkAAn
hzrj6w9oNMn2FRUk/9jjltip9O/EovGC5f8VilgdTRi0juC518wAxdnLFOExMz5roWKzBX4ow6Xd
pixpF5I5kjsXqcjBAYE4/tDBzKNG1drVk5U+o4LcHsEIJ4Q/FlxFAjpXl6HHTS1wrK11T0AiKZBP
gjVVGKiBqSNb54d8hXDKgWf4lErQg8bDpbqX5TIIKSrcQemRMDDZjiOLB8lc7AubMJpF1AParcnr
ZkGiMd6OeEN31gADhrycOpeyMSG9fUKFu+RC4ocBs+lCwCA/8JXrD71ZTIZH1Dd/MoQKry5ZQ+xo
nx4Yyxscc2RovFLQI2p6dIfwYHaHdJhnu44bn8N/YNLYKm8ALBNqaomr5ZbwwEy+eYtUIYu2efEy
dVsM17sZy9URy05s1CslsEz09UVbTHQsiK12U9tCqYAhFVL2Vjk5BmiAXFnlywbniNiqdzuaoGAv
31B3+ZyAbfGRaWkmZWcbNl78JO99KNRnp+qDqd2OLSAUBmlBYl1ZQokfVQtpj1EnFGGF1KzgAn1/
rOew+Ka+kFcyOzjl5K/LKTQO+dJfgiF88Ba1ngFz1VLbSOlZHndecuryYituHnwXtItmvqiV1LtO
2sYeBus38FXU3phKeeF47em6lddoZ9TcKB9y1fclkJxrhMK0++zsOT6H9YE8hG8WP4jYa8BEkCCL
OP0XCHx9Q/xSspHosWDT8IYFxG8VtA1VcORLIvRpLhSTYIhVqrRJ9gJeTgof8mKEydTR22vIzPRT
rZ2StwO5kYRWvBppq3cXMUUdc6y/kx4kCzHqX7cvJrpWH7OmkRxTB4x7lFYxExACVYhmxaRx70Bh
34poVC86gBIrcfWpxp59P7/9DIzSP9PTVhep1p+M3KMW6V8d+p1zNrs44oFyUQRLbp0Az55w7rfd
xvMYwWA4RH1muwG6Za/gAP36qXs9/PESgvlLvdrg8LkeE4ilDXRfBMU/rK11bFgABwTB1x7GTGWR
fCs9Tzi8RBCa7NMo2Upt6STo6Y1fr4eNL8s9VcxadAy4Y9f2KjVKuKAb4Ds4c1Grgg6uK3/XFn9M
7EvmY99zNzyLFsYGyrbduZ8LMfY3fiaDX4GXs1xIsQmTrdJtN7Ew4xFOZ9NKsO2E08kgzrx1Aeiv
sPUju+Gf0SBjjixegU+MzrmjVqD5CAoDyYJ5N0oWc/laAIuCvrgbCJq8q6jmL/a+L8YjmxAMroDM
yoKAxMDyu/IAaDWLNTrQctMOdMi+dw6wRpDYQy5T4yhoa00wH0imjVIU+JuIyXK3M15AHbXCXdjs
G5I2H+1Ji8DjaQZuDCNUCbBnx99OMRKe/iXeukJuBD/gH2F+3SJxtM16oI0Z2gWAJw8f+fMOtbj+
n348onIbS0i7PtYcIARvoeV6Ry7AqAamEAs3Ber+cEL7j+caMke2F38xsOZZvkAqWo+AGeTPSVT5
7MNIva3FWONV+nyNGBHi7ot9d0I+viCmSML+TLhRrpBBDl0HLkvCR+qwEVbRbbPHdaneyp6i/5J1
bWsDEfDUaHAwpZSW/acWIar847DPb58Uay1HYkDzSmgYekepm/fJ4GuaGHfitW2BZu79h69Cn6lM
Z22ARX66Yt3zv+LcVey58IvAxxzssgZoOE1ljZJWjz49pwKjHQ4GC+kabAFLJ1LlcGn5gj2tRlM6
fnXceOg5luELcJ9z4wTUkplUK+l6kMnXs18FN5yYfze9r/QbDuh5K/MIn/oDYqCscf09/ML71R80
nG3dXQTgVj5qM2S+aTWeGuF7Rhh7tmrkvCzLfL/NyefcEzOdcebhBbd0f/69njCKiBGhh0uaKzAi
A4raWLy1f8LXqUYSPlawhXjOZu1ClZ4V2IkaYgYsz9y2LktWQMMg9R0+0WNziVKo5xfOZU9HrC4U
fYgBOCkZ28lw4yCepl7tfpacMsPSwZV2ySIjmxGvL+P/GD+pTLyTx17jJ1ZxINN1eUgZuqvDILQv
A0tyBjNDZbBiibKqm3rG2T6/g9d2sooWNnJlrppCQjWfvD64fEPLQN9dQ9kRIrcuP3CrJChnzOFZ
GOcEJOE6/t2dqjNVMPIw8ebI1RG7I+e//BXP4KIgi5w2KQRLS1OT0RCpN/BJhTz6fx8PJoa0GBOx
MbzNegUbaDcCtHU/f8pMeOJFF6czyytQKyUqj2OMcgX+VSY09PbKjk0ZK4COafCcY/XNqaOUtugi
CSX3cKhylByf++fgzjX1ZQQN3+7waSLSXF/QBx3ef80JGblvQKdYG4gfNbmq9oIf/+OqdDAxLVZV
WbCpRZ3R0zqkHcbU9uBh5rPXoRFLZNafFuu6uYzF8ecqw4xGoufCmuHa+AJYwa3o3kM5/gDotc2l
D/01mvulV59dTLdlQv3GR6aQDUKxiCMxlH99FJD6XEy1ALNY7RGPaEKBty0iSNB98avU2TwdKuI9
n27gthTmhsmhl2+e99W4v4eSLzxhwUCBdyJZ8iQ0C8X+ja5oEmF5VCpLgjJZJbvoXWe9FiNlfPNS
mOQLmt65Idsku3KYC+tBKKUl/OSh2QlRHSSQDYup/i47lJfLAx9r0xWmBETPLD2GY/zz3X1+i/nC
jhEXW3DS/w0R3m5+DpgXiKPcNoIHVNXzxncNDAnMgHEws9ezuzdMpEY6jEQRHwVhW+g45wqo+KhR
7QpIy3Ykb1vy0YHM/DiU91YJmdGK5xZHatFB4vAZJeGvp329XOXBNRXlQNfENsh1LMnLK8AEkFhu
hUWpxKatIhJi1OmUcD8VNUDhhJ6MebXj8CZt0s2dUk3qX4Ke+Ybz5YioZjVFGaRTTIIdGmKheuai
qpmUwfotR/lpyGc/QM6eZLCratVuaeyxlLwWWQTHdN3OSKBFP+OmFYZDwC9eCdU0qkN2LgNzPInG
7G+EcwMuFn/U6Ah3zjtYz8cPqkqI1g8RCWsRNskYtL+zxWWxQj5STYYJzRkR3pNTb9IbiO9NMiVP
daLIZ07WfDJ9ffEXejIZEvNHuPrYuwqOtNh9J106wlxQ3WAC+9KoNd57NiyBFdfuanwORtJhfgM6
4by1SRJfnjPaUYdDANgSoVGYzSMLwrYMIqg++EN04u65lPiCiXXsUrijoFmbP+Oi6WKbJbUW/dV+
BBW6TuPAlyP6YH2agEXA1xGvvzvnuzQZyBh1MH1u8ZE+mLvYBPxfVb96UiHY9bO0lCzZRBkDXJul
ak3+w9IkI5XZn3TzWxsw+4cbEyy8hRC6hOEJsSi0sIkOexI+9yVD/TbsOjV8PYPfgZ3/Wer3WB4c
DpHejLO5JRVcwzNyZNGxC1bdI+JGYdhnsvBwzmD80i3KUh3CSmRCDsn/TFfzM+3Cu7j6DN24dk8I
/Pjl0Vwfmo07+wKBBJufz9d65DBs9P3CvoOBWBWR+BrCmWQ2bQQ+LnsTw6pmvV1qJBD12XFX38xg
BC8Lq0fqtoGAb5Cb8ZTIlL9Xcb03CMBUOE06nesRXFv4fco8y3j9HUbH5pVWtfoGf2B0jwpGZkG1
jox/cRDJZenq6ukvqWOHNSarmurKu7p7XBZRRK1eyFHInykRZ+HFKz6DX04rW7e+/uvQWDtZVaJ3
KVtG5wMNnEMdhXkLLpReNbvtJndxf7G53EMUrUWV4rXCgOMXV8S716yDPjZKhVAAl0XkHY+ijyZ/
sVCsHxMbkv8tZkB5qRx4ttwLLYucJ7iBTLkF/Oz2B97eW0lpnMwI4k8oNu4THCZTQWNxhGb1OKdU
41AFPpq7w9e/n2O6a8hliv30aLeYaR3+FfWUsb8L4siPzkdahnqwvzVx1Lc8CMv/KO6rPCcYx3x1
TU+w1CdLJY2of/1PKsQXJw1KUv9ZiQ00fK4rBkv3/WF1owd0eXsOEfkBFSbjP7uPhFxsqpxm9AK1
zc2+zLcNe3moVxERXipRJfBd3f2XAPFMPEYIksRshpJ/+izo2IBtRYyH974vZKqn1y889m2B02Gj
Q3ZA0kDxaiNLIO0mtbu0/nQZ8PLNrX/iXQrWPLdf+R5Lsq7j9GJ2+fGEq7SHRJJcP/h6o6P317nt
yn6osv8DmY2giOZWgA5brxIWM2FgUTXnMvajHZzYpgjjk+Apy2pjLYUI28axgZDkGpyl9lZf1QF5
cA2X+U07T1gliO2p0b//cP6FXbpCCW8p1e97+0C1UcPTAkCW2Wbtk5iQU6kW86oPkIC5Gijqn6wH
jARA1mhTPZkc30hM1e3lUAA/SQgLHwcRzEadJjmYDS47ekqLqEKmgL6+YDvCrB7yxNf2olQ5DBe4
VOiqFfbKEeuL/RjR4D+y3o0txhOMt+dEzG4mwydcV6UH69J5PUGzS3dNDb9gIN7IXkfrq3Bhex1k
kyDnTGGfeAiLy6MuYHTkArkcGrtpDH1quKaxwr/6N2K7VRMw65OwZfMiDHn5Q3lWMNgbiPk99Hw8
F5dqyufyDwJXA3Wnd+BySF4rRKCodUWbx1wrh52WMSNSQ4kBz4soKliEdXrkYiTFt7qsBL3ijaw4
hw0eH3uV4NXZ0LOCK9E5Vnz/GEzvoaraNzBRMxhNYw/t1oR5lLcX0UpqhwENx7mYvKMDIVZfDYT1
+T8fy0Wqcj6uiqxvCBD1ZUY+yGflsscasl2Wh/fZVO5Pc8MzuKMxLHhvFjiU+LcBCg5aM9llvO4I
T+q0kuwZ3hVHvzeF1G5A4Qz2M7aUPTMnVK+kHq4KnvZEbAESaDm9enqPa+WYNtkA19Jp03LseSS8
/KM2czylAqhwrGRSfJPmDjQqquO5JuXgXbsRh5FKIgcVmZ0kZt7kdCHwhe+OWzkSznLJfvoIh5Zk
25RLCGytGyt57WBa/yD79Dlcwk/hqkBzjU4r80qqE0uznM5BOQ71clUOEGz5bN64fxInadyzMOvO
pqAGIwwaFzc7xyna5ryDACoA6e4HcLJoHCIQ9PgLq7GVxo5WRDjcY53t8lkw+a0j2BvwQu6S/oX8
E4UQiRIpL0s+zh8oTDIM1s1PP9T4OaV9RP9iOyOOUAT+ITuZIY0aUV44ubFpTXq1fOlN2nOa7MeB
cs+ISD0yrkjCKsNB8TIgjqB+sif6Y7KF7cMpCJfJtUeC0kk5HVXSdEHlkLTAoazoOU76LUfY7FQg
783p2CTKSQGBgMPyBf1Aj5gGfJbyoyBj1gJk5hBO/sAgsa976KhEi88QuRJZ4PfZ11+VivAarL+a
Xt2c2lZFUAISBkqJJbji5sHSZuAILPoIps2KG2OGIw2SKtxYvW/FSMhNHLrFgenoEIXYBEZNtcTN
0dvP6VY1jupp8ne7YUoXoiPuDrweMBIUNM8qNBuHxuQCYkZQZrpqLqNd4GLdLGLoF8e8+TvoOKbl
bw2SnWqEkmjZfEm1aWrb7p/X2IwgILigkJ5QDFmrysZdchZbXKoUKhkNZYtRis/9ptk8MsqkRhn2
3CZoBEo/8fPxEGsGcf+T4sWAYVq3d82FLcEC3/CNmpRF3xQCN+3EDwFOBKkyVl7SoQD2TxtlQgK3
aF23UmkTcMhGXtzBOVcjlWkjL3P5eCUewR040yB9G9hrxWr5/AFLuQgT1bhbzvAk+7j12WK8SYhI
QvPq4pJt+WgiPSm0QRC04Lj5MzyeBzDH4Irc5sxdOjoiUNx7xktLIGdpJWpZGpTJeswdkOiwJLXC
zUhgK6WufIqOjAoXYtYsjeo1vWC53/w0jU5IHKVYZwpJRfJ2XQiQuDFjI2W5TzfafuqBPjfwE+Ve
DPVUzTnlekGkVCFwSPYtGmXfh/9/p3T4zKZ3aeqibW3M9fx12Qa/orj8ICKVuSvJI+Ys7fymBQE/
HpDVfgGjrZE3CjlV/85AOjyVohN9qKTuDiEar+s+UAxP3HMa1wr9fv68c6YCxdxiOvihWmaSTINl
Hh1I4Ty4FxCxwyuCDgpCAiA0o42iS5pD/GeUyO3ICLTdcNV5a8xE7GSlkObxKobh/M9qn2KgacNY
KtSzN3vXBpLyA1TFAISkU/ImbeO9jke9AaC76Vn1wOGcc2kN1ZwUdIeN8cCCGSazOO4hvPAkwVTD
WzJfm4rxSx9daV/XsOv09gyWq482OXaOgZXe99xbZ3VLjPVwN4/Lt5DKp/06MhjG2X787iOeeNGH
RqhXjPYOMwwCiW8zIl9NXC8dNVRLVeEELUC1lO/8SpRl4uYOGTF43lLaaLuq+hO2lDPtXKX5t2st
7Ch83cPUKqeD3fWmwyryE3e1dHnYBwM62v+4yxwIgIxgqIwtRZvtUvY/LYTErfN6Mh/Gti/ayrPe
/tiWwHcePi6wd+XXAHz7mH8DBFZpSewrPSkN9gBqEe0+GVb29PEuBjl9owMLYF5HbYOAUSL15jaY
Q+c4yHeMFJLqrQQFphfkTNn3xOTcb+KxkmjihEpxYvVvY2OU55dpM63T5Wl5VYsdg2YWrNnds35u
p8kRd9UA/DfQKS5gDYWfTnQ/WZKzG+O7ckypK2rZrJ5n1yY80CQlsSMjFKpbq8dfrojn3W+Ksqtg
W99FAG3vvrgWngpD1EDPvcVq1k6I6bsSeEhkINStmuWTZarx725y+sw31iomeWiwXpxrMkqaCX5G
opVV6CxwqeeAcT5gE6nsmO3RGwbHJYJInMCF8jhsjj8PMpYW+e5NUpTG9+uDeI8xVHqozX/HqfLT
nZOYToLLrIlNT/t4WEwBtYkeJShiJXPADIVoPoIh1M8JnrZfULObDdsbfTJzI9MCBvo8SnKWjWi5
z2qkiHEV7lCpKCxL6HVEA2xmAEhiYR1UYx9/FTGLuIqD+bspN0XZijf7SMD09W1p2dMZqClqN/hO
Dn+nc7vUBsIFwUGvNiXAmJMk74dsYM37vQW+Ls1f4/3iHKTm79dkWQ/7Cewswn+mIklzB4N66sb0
1iNs3SXjTiPvzTGy5eQJzH4/uUufPNn3gYTHVZufZk2LkETT3TDvelFFNVlaFobQpA31LLUt8yUg
d0o34qpS3NQ2Szih/bmjEKb1khLUdwJ9oGaVpNlnMbiwNW4NpCGwQQFb+Ew0rOD7vOo4AyCR/aL4
MO1Ix7uVe0FCNooxuYqNeVMSWVohE8tGOFYVYX0+SL7vKeI16AydlyHeT0reTBZcClsegG3LYrar
QAo7LMTThBZsNKY78M2qyJY5dddnUbZCmVlGJrqOok4jiKEFDF8GhL3Ojy1zqOi0Xc8TLsHZjcs9
I/u+ePfhBXKgFdHGm2WRfAg4mRvxVd1sqYnNlB2v9rwF4PVbjh1KVdy/78IDEg3V9Sdc4YyYYxlN
1x3Gt9wKHxIp7p0KfzRA0qXbS+TS6wZVvw0PgRA4Rosy/vZjz0sNTRBbZdh1xRzx6oxR7qBlpgw1
rk5nKU9lC3oN/G59nVbFDmLrZY67NoX0DG+m3ncelhGDOsgRB4rxLA/Wpc3Q+/hbuGz+UQo43HJa
sysO2eokGLi8cDqmrl9wuXIRrruZS31ApWm4soTQjKhY3vUFBhppIwug287iecMKqKuaRbYZwcKO
ORFEAMtcPK0scIsuG+g2LNw3B5UxzWxqdvcQ5GqB4mTg8or5IpKfDdSvJSH/XGyeO6/F6NzCvokT
qCLjZqDX1zuoGwD+fFCjLvXKwXUMNJVcEY70YLO6Ohi2UDFj2saynRv3nbpTCMW8kDX+Ev0acKAN
cOOgcAVmMSxjiYpVxYmRwyZyiC0XXcstEIFL0q/3LrMEX7I2Q035SXju1V7F3jHsvMNmtC4dJhVH
D6EF6UQRqC8wKrOrGWHfIj3eJ4Mdk0oYEwGVo3H8lm4rIGs5OgLgiJlbecyttM1zKZV3hj2gQYOQ
BRoBCJBwGT5Ueler2fedAYrARIzLk/kcGR0XtO/JA+Cjs+rWq/fHYlRo7NCAa3sjH9KDjO+yxrwc
TWpTBW+5eH7nbo0ozjJxgsrvHMc5tcr8SaCsxqnNoJ3yVv6tnt01+ekl8K/dTOX1Sn3u2+/6eB6B
FcZjIa0HOm5Z8s8QoyGp5TdFI0hfn+VeHQZ0MwLI29ATeSxB8JkJv+eK2CPMlWrwCyDBFTbgf7/1
wb6sZHREe2zN9jLuNdAPKwXQHjcphXK9cAScomT99dux1QiMoohmRnxbyjDlEX0aVNMHAl1r+nJP
4TGxcDpC3z92lS6Eu+Els2ajbvxRrGlc1QA/+/ooqE1oNl2vsAdkSnB9DrsViTLE8f4Igv0ShYaV
6/I1dx7Z0F1Ld6v9OI5miSdgBupzq+B7bOoYjAMMY28b3RXKf8EoueQUdjC6OQy53/Zdj1VqfpP9
PVx9felNBqpsZwLFCpFCJu7LbTiz2xRYUYQoz5PFh+Z2pdEgxDCBejMPG5Rit74r4Sj7QuMV1jT0
4iS1C+iGy8mukcwxoPQUCsdo9frv25qnH3rwCdGQA1G2GelXzTn5X27Q7XfenEXDALR7lag71cdO
hVWapjXDRFQyXRFlyibQAdc7b5JWLBjxjrr8SwkaNCrsTQAy53OmnJGuIM8tLhv5dbPdwDIlpyzl
D1/vfv8Xryks7MxZ2i+Lr/7kwOp8UolHdBUC0A66JWBCVdtk4iybV18yUHWpYfGj/dreAD6YFpk0
N9toZybeNQsapkn0yDR1Ai/NcjyvHfJn/RryCS17r/TTADqy+By0OSFyT7xQY6JB7jagPrxwfHsj
OOtLU9UhAzzjuN7UKeLsQHcqCEis8w8a3RXYsUerrdL1mNsam7ZZsyRam4EBKVYrATdG93V6imCz
jC7uID1Eichu0mVml8Yy6Uh4HV5E3nooiZ4pmowOmkWCOPu+Xg8pvRdTHKu5aI8wE1+KsDPv0xiA
guSpU5cf9N3T9hh+2D9ZeMzOzcc+YDTpVsPEwyg2JW+H7H9zAjQI3AkVbDroO+HBaLXpct2nP0Z1
CFCPWO9i4K8uRxQd6bdX5hOMnpgvZ+hv3d7fCB2G/V4ff+VCC17seEeK98rtpLdr7CQsTOCem8e/
cASsqv/0Ki6QNiWl2AKMQv5eMTutoBUJdiqwSV5so2goVzn5grxNrschB7vNj2Nlkhr/7GCq0LtY
A9wvtpRaRR9DYlpGclft+ejCIXSIl5JpiPgPIx5B1ZlIHHcvz/J5jv/UymBWMsulHOhUAtu/EEAU
4ai4hqvphmSL3Wk9CWTNBZFG5VxFY7VzkL/OCZgRRPkRboY5fcu5T1LSxdszgsAXsqw9DFyyGLoz
DU6zoK1O/tZw5O8sE8zKTB3PvHz6iJ6FdG4YwokjqmIvvkyxBnlmB+P1q4H66I1XCDXu6hGY0LbY
GO3yw5yHCbueamyTic408d/TSnlcMFRHQ6ugDydqysvfTBCJlDxEUdtsBvS8ythjK9DQrSuWXNgi
fPtW4x14ha8KkywHvIV59Xd8FNuPhnyZRsyhydB6mObOdU3T8qOpPGHIMAt8Md9D5aCKq24NN8QE
rON4zRpGvpCiX0IqFTRXdITQPhpo+2EvN3stXF4wO9T9Ucalziv1yhQtxgm5EbxmUjnoz5djn0GE
c90YblWv4/3fZqejt4W3HHp2KegGl0+OgJR4ZlNUAeccciPsWniPERLOvXAnpJoaxfZ3N8aO2BNR
+vkzajUq3xly2tpilrJoRmdP+mdjLCbIT6/mQC0fO76BWGOghcSoy6r6JLXIM5k6P+ImN0gbv17f
A+HwH/+dGnXztNQ+RGVyAYNniGX3YEsLhTcuYy9hmSp/FOzdgxdjBxEFaOeAcDe0Pb5LMMMK6k+R
SO8h6Jzc0lBiYNjESFer+kwPX2AP49DQaocjsM8DLebM+TwCnCff1t/ud7VVVi5uM8eXHRe2GPzb
nB4LByVwbxthS7sMTjJHH7042TPxEw6YyeglAhJQ9LxeSwd0uhlNMPBXdc5+RKsCR3Uo/Ou2tfZu
FvQDynDRUe+F9AEfJ4b3JILGyS2LUw7A8IyGTUS+v6RBCnEhhaEs/Tqh83CbvRt/Uc+Gn+1K+riR
irNGlaqZLnL7BZRbkl9GeZy/HDn6zOkb8Oby2+CE1ajKMBpCg7YAhWpzBLK2iY63pjYDAUYSXCNV
Fn2kBSHp/Bb+q9joT3pa+S/W8PiTRHwgHGbPzRK60mYefX4MBDfTrDch1EhW8L2tl+Y6R5gtHhOE
BIO2VlSa+da6K1SpYaC3kzqIBsKWHKjWVrtohUkoc0zF+ZowOudLi5PjLLDycZjDut1S3bwDJXpx
6Tvv3cywH3gl4i15VDujaRXitjl7FWU3kvJkGsCtz+MjM05dMS7Cx7W0fCD40bfpEzVSMmF7CwiI
P4qPCcpctBZ/l6fFCxtD71J2tShTQzybtcOnDS8jx7as3G9asoS9qm68iGQuEbDHq3Cl2wfjIx4f
oXemPWo0kVl6wvHzIvn0tawP/bJhdpFsk5A8+Au29U1bw5HilWLDmUzeMKso187ibntUQYE21N1W
XczN5soSW1L0Ra+7H07ww623Q8iU8xv0l9sc+ouH7SbvgrSLESudv5Pey18q350mIyn1dlnYLpJF
qVr0kUwlJ8SSxPCFFWjK4nvxSgTmuJL7ZHmm/BcO2Iu9EiyC9VVAVymPwlEqy/QNWnldYe2iLaha
K+vzmaNfRwPp7sPBlscycLdfESz56cZHgsRBS65DmRHQG5xj4SdtzAKdZeAXg/sazjwVtYnCyRIs
5N/TmaYuUhXpTuvZXkU9CKrSzKyoI8J6LGvzz1msVU5LIAARueBREgXVDEeKpODR866wyR96+DDW
uaxXe/kkwQcLE7YPby+jPCB4VCZPab65oOAojDnkRt5wHyYlAPkCRBJaL4LMLn1m8s734qoT1Msz
7PxgdjoMPBZ1QgjZkIjUwd/jn5ciNr0ph93SuSYS95eNaR+YBRX9FAaCCP/CEMemP73mq6mROX+C
mu1VECn7lIFcVWjj+fcIk+z84PGfvUGJt8heJSXeQNmrT2HsqmVpZ7SpAti2CQPkR3sQ7JUxN+ly
JzkisnkyFYdzd/EaZKTbUeAxgokh3NfShxYTAwK5K5H5YOeA3er7bE/JUBmrPD+Rc3pgsTjMJP03
wM450xdIkX71o+aytkVNy4G1D3jJP3MsmPCS440N1VA31zcYV1PnFdhvmrQcrlMTiqIsr9jEwfDF
7Vow2x3iOx9psvxRPyYmfMHqoo778buThyVyVlm8sDfo/p6HPjb3zfHbK7Mamdc8lBRaIvqQwQ6C
VQBA0FHry6tPjQTjJf+4tqmPelZ1j9B1eQAMlw89WEsnslLELbq4X55942E1UFD7y0VtJayaE8PN
5zBaRxNUQ0fmvU7b2k+OMVv3O14HyYwtSUZ7CLL3VhhYfz2kJBytEizFy+ojQ/1mQwlbSWWTBW1d
zV91xD/1JUpDJuCDaisglJadNzKacMZSy1+Z/xRv2kBfhfJajujDLooH/W/kPtxuVIw9AjSsHFO8
JT7XBA8O++iTTHmgPH3GhbrIhXKWkHS7xpBiJma+Nb7RhDb1NdKwCmCb5TaJF/hbhfZ/DyhirD5r
apMwyev6sVqumQRder9kv8DLyFq40HF6QDc0xovAVCVqgILJDciBCJHRN8V5DtW3/Q/rfQCnhTo7
Wf/G6hDIV1be4hUKMpv1xXwaiozBrL/7RNKCpege01Ot+FzH0IR8BKA3Z+/PjFTpxcsNip6kgYil
WzhZ+xkNFe5Yg1Bzq9PDhBBCwn6C8r64UoyJTsKG4qXkHjcee8ez0hi35CpQTZetszWMJDftQX5b
1lqtvm5mDqOKKroqySx+Yl++dHQEWiSmR3KuGm95nGlrs/YhDYSeSI+pw7YTXJc8iStdOCKV+2oC
lDG3WUbkncRm/ER6i3u2xPxqwOQ0cXiCCF2hdCamoXFig4Gji1dxrtbEFjGkBM9MRihvyvaSuqX9
gQW9Dtvp91yo1UuUuaCFiM2CDeumtvaTLzzMDs38RY+V3EPgWVpvOR7nRbSF+J50352ijF5ejTzE
/RvMz+/YBj4m8og6m4nlgPaSesXcPMwDodUdimJxKcI16Zf5AqMHmOZh6R5SfZC9KpPLpOZCj0Ha
RbnPP8b6vSvr1d7taHtK++Yg3miEjusCp0uF1h3sXWBx5/+NlSgz+2qQPJ3dDqfU8eSr8KYWZk4z
2es3XekoidMzINHXJyacEIQSCrJM/Se3SNF+vd68EKM7Vp62dNr1+QKLGLIgM0F+UAFh5U7WuJDv
6BmMU7YPnGzwiKNOPsI/A0wqLhuEjD4YrQONHSctYXwnfqrscYgYBs/nB9QYb20wEOCwK/xXzLU5
md/0f2FRh8n9fret+fLjS0xVYPRHGsdQWCDw43TE6B5p4r66xS8GhoxM6NasFBPbptZjaU4Y09x1
uoQdBp8v/wv0sq9NKIY47A+cE3Xns/UxBwWbON+5aGJPk5j5Qe+Dgmtu8RYYtmxXAs4dN/jACAHO
rEtJ4wmf75Ke2945vUmP0HHEssp82c02d0LkLtbZYfOg6RC1p4/X056wEQd/h62Vj43k/YkO8YDp
SjD7uBL05BrWKb+tp4abypYAm4wT1PCAU4phq9uSAU1k6ELNmcwHndjwUfRMtDwnphD1pm+yqmp0
17bLlY81u/82d68OLnxDJhKQ6ZZ/aTL4AJaO2Ehb5SjVULaLZ4i2G0o8ezhSiU0fK3eqHUNrDzQm
YQh5f/H7yS8ZBkzKNtGN1YMvodtnHE9ygIcgnHl2N+LUwuHU95aIutVj+MnvxgozJNDASP1jKjSA
J1sLJ4rzYboZ1dsvoiATVDBTAkNJalk1xvm/mFl/jySY4E+hSEmzY/NgwwPLcfG5JTPk55eP8lVy
z2dbJhkc1wDqUps+glOK3bP1/pNRW/qXVZ6n0liQzGCUJCJPuMWdheluWLcFhd9eVjnV4eRMEK2+
CK3cNpnISVqBSkbd7LWDB0Gd3w/zmAoCL3jvYNlK9FoNNa6kYWDsjPFVk6q4mVuCmnWsDAcOEQrq
QvTjLQmotYdn4sa2DcqAmhiy63dIwrMqfSTPwSghFmWqTtgll78mJ+3L7/EkeB4DFxIIugaq+9Pd
wozVFlwTYMyeVF62gbrhErm71IRdApT+SRdPOT4s1FNZwp2xEBf1SC8FQEoXURP/E0ufZdE9L5Xg
peJnqrXGlHDH79XxRvlK8DGBSz6qv7NGSLMqrOgR3YlRgns8XL5oNx98cV5qAd2kWTptYFfCllmX
ddUWqm9DaF30CJAEeC4Y877TCaJtxCaUX1D+FzK7eT5ZzNkpekLAW3a6ZKHxTPNCSniPa1OTAvPM
xw/gnacOMMkE5qNQGTu8pcGevsb0WqCyysWPIk3ry/+0MyUdwV5oqth5MZAw+60AmKjW0F8IkcrD
jQR/z+tRiz5wPHa3taFqO4Q/E9ck6wLd8NKNp9OpBh06roCyM2kfjPfsCEK2Zk51dOv4QgJqiJFp
z+LRNBSsVyssZBVgCJrxfXmVRGuYdNt2E+wcLFIfC6WYkiRTEwjm59e8HS7Ku7ufp/4FBASG1+To
m0jOAgjkc5Tt431zYXLvkwaY6YmHScRqRvuUZqe/FAMjqWFqEs+i6eS4EhrO+lyE+KMiTX/Fso2n
LKOwOoQZnXLhertW2SIThxBDr3ucPLgGMXqFt7IvqKVSFzaps6Ua9Vc3gBYW0IEsf/btdycd+oi9
n37WcuGmZzfAYqShLNPaI7Ca+4iICTaYXX/RjSNFJiwMhYxx7l3exLGXP0E+/8OGV/thp7FY0H2t
ALC6JiEMVKYCaAK6UmWgS4dorX7IW1pNqmmKzgjPBGw6UN2Z6RROkp2M63lw/Kj4r1RftgP952LG
/KVXz4OSDqVle13P296Qbapt0lqWKqjNwUzf7JjAq/N0OsyN2I9Ecy5sIebKCsRvgXL3Y78J+62G
r2c5mXVW7hpg6IoSdc2jAA/jU9YaxfwLTz362Et+Enkd+J/caZ6URCer+3I57TE3NLXJO7MY1Oxa
BzjyS/SD7NqmpUellpXPD3DIi33qjls3Dchc35Jas8E+rYL07l7qumLbGBbe/VbrLP6RU7xcVpFb
nXF+hLU4EgRvjGfpZbPSIhbAOaEUnib60zpXIJqAibPcL+MhV/bz0tLHvSZo0yz8yRTuazia3WVn
4VPTmAD4e7hu4jRt2K7mOvb9wH0IFPdgQe/FORreLqHuWXQ1ZTW0thXA9Sx9xYm7I1KW+Z4r5Y4v
z97XSq7fsimj4mQShhiUkWjI00O7q1Fafr1egcprgRpoTdk7zUg6Xd42PnD2YZYWx8cEqfJZH00z
hTLJ+2eZ0Bbl4U7NTsA24tYRYqP4wBStZwXbsQe3gqDdxpVLr57QZF3PV6QfLlqEWoiV0oZMPzpn
f1SBO030UPodUaOzbzQfmIC5J0aUWcNFqNumhkJw/6yKfT02cq6yAQJKXCZc+PYYL3Eydbkt3Euj
8pbZkx04ZX372aY9B/b/UcjTNzM7Y/8MjzTT460lKZzJGj76wtQg2PBF71APT8tVlguvsSDrHDIH
/rnaoKD5teJSHBGzcYp0MbpWMj+GTw2g+csslLTUPE9H5HywlQRWqnvEUKLrirRJ7N2VrJjPPCRB
ZELW+Vyib0VWH7Nv6sAbbxpf1sNqMeBDh3rMXWyabRpfbYs7Re+atiEqPRrPji1Be92IZqZ/6j/6
oMa3YcR4ll5KHoDgmdR6aCNFyrFsZHJhRcio1lpbHAl8RN9p8VNVQDjAX/iuaY2msZW5Dzf8hnaX
6yExGbGBI2DRVMuOwXvenASyJ/T8mIzEy9hNjcKwbyNPosnRWvuCd0LeJtZC1rc5o5TABA2+WtFv
owQxEaEL0wZAToscVm7qeqe9SAPfRsIn5fQN/SB3QrUVrosS7gUv1HueMbCHny0yRmPAGOqo6PcT
zK5csiDnYJsUwlBRndHTSVh19URpxVNGDISKUnmj7MbJCSyXbMVACzKxfX5a6Ko0g1vVPoSA04nO
9vwKCPkQporaBmgjAeTsC1xGNwN/3BrpX1nanQh4IM5ykjFZ0nXc0F4sU07h00nPhsBWM0qG6G4J
HRE2srPeAuAAT6X0fEQLfbzpYQiTLolyaNqklkV6vopY/9f/QNJLTkNUyf9BPTcd/PTrbYDwc+6x
Q64X2yl75Pyek4+F2d68biUtb6D7jFJPItSDr7+PK45duPER6CQrGumgw4hktlXaWcKAOcj0MVmI
4XWf3W/OFBnkleBs5DOgY/BeLSx7SPktIJQYcBpEmdjwASNF6VKcWy4acruyEeOUr4Mp1P4yS+2e
MJ9mPP44dYNdTzpjlAJRLyOC0e47ecsFPY++LghEO1okEgc5Cc995oQAvIz22s7FJr7Nyfa7B6sq
DRFhPbqOQxO7wgiJB7pBD0CFZbk5cdLv4HPRlcVBl6EJO7MnlcTatfFDGuj7LZg4369TXtlS9Kgx
SqiKH54WPlvrnrbllaCn/nvd7ErZNTxL2/1sxz8k8hxxIekoRNm6QCUgISw37mi/GyUB3IJaE2/w
M7XwN8lCnwm9P1/Yo53rFAk0B9KQ7NX8WKizlO6I6tAmdtpIczfi5rYLVOG8M0OjcTOfMKqgtOqb
oqRqIJzHuxjv93ODJ+7wg97kU089DQeBrWxi/TutpW4FpfLW5OSPjkcMhzVHsk0fqv0q/K//yv9Q
08UszZkT/RH6XHc5LrIFQVpf8DKcPhImMWnjEVHQweNP/bX06HDp7dzl14Q6DBg5T3pxCX21anmJ
IYCborht2If3XPHeNKhKBUVx84t9ruUqGjbvexWStsLo3nfph2atyEuJmdYElU8t+ojui7JGWReY
sRkut8ZEK5nSflbZm81QxBJLhrUzaqnx0MXzTsWWWiL4vAsbXXUBcrBgdb07LvscODw+YetOmN4n
UCFLMFqhgf5KwwOusag4WN7lAvlzQ4hk7qc3yN41Cx3HDdyOOpPbqIF48kTghvtvUvUeAvFMgA+j
XiSEXhpInZ2hWrkJ5VGv8LGbY3Dcf3JX7Pyfr1QimIZhCEA7Y3ZY5qQCX25m7AALzmXgzXGETpQz
ripcDz99ObQpgUMn+/yF5t4E3eIXtqtXClSJ8Xkyi7UTGoc5YU2QA1XHnUOBb1L+vquxrmp5ZVPb
P375iW5uUMr7fuwrAUvWw4NgWOBDQwG8yacLCS+28ruN0vXHjB5civ6JGTUlecKgZbCuws9gKNcS
uIArS5mW6a6DZfecjhv4SdW3hgnAzkzmjJixjbNXRsDJ1q58Lzb0TDOc21fvZCam7eSeNwsuP7hF
QZcZcjD0isJQp5beJAQeWQWgyNiLOGwvdXJtmyYGVF/sNQrMkbm/Mi/Nj4DY8JxknSj7wnSF6Rrk
FiG+qRvltvJKVdf/Kh/zzLWsJZxzeFQjkY/jrUQ9Aguaz7skf6Lcq0p5e1IuYNBBPToa3IyNdu1F
dF1WWNLpYpowmSDNyT+o6CBz+FeRFHiYN1vo5o6lctJMdaoQdimAGqxwU9fQeBayRAtpFaECwwMT
nwsY+KBNUcpbQRgRTRtvbo9GnZV5mz5E9j/oUCdYfpIJZbHllpGEQe4STBAU5lQu9p/yoBjSAdkG
fDkPkvACz1sy5LIfEjb1KxqVrVM+ejuJRYlm+8ISaRUMMrZDernUKCV+aN9dDMqNzuEFBwOM7tXZ
UvocVfWx2FP74kNWtapBO+DUl5sqEv2amzWUjTFFoejoe0+3ztcixqJao5PueCn9TjI8BiCYsMlJ
xU+KbyOvsEDL5C6hCkMkx8baT7v0G/oUQs76Y6wWUKeV89ThNdqz6sYvUCVfgeUg43Cn8okq740g
zPXquJCO+pIOH/Mf9EcdwFPdAMn3ujb3Sb8neUEdbiaB2x4KAn8lB6wPnPxDEjJa0xGBPXvkxd4k
TyWpGMDvZ8XXR9SQNWemR1tWKWZZfIHOM1iCB5sBlgYBLI4tZG2rpn9/zSFxYhQvS3uesNWC3+MM
hlzZbwbzJs8L0SfMw6sm2aWp0JjZnVSSfeNog3NSDqst3AZuL4QMQZIsT1iBmL2lAZnzD9C0E/1k
ehDuG9N5Ci91XGTHyJs156AiQSCcgDqRzY6mHs51abNTtBmwJHKDNcxQAeDTC0NP/iLlwXLOLos9
DZwr6oOiR1yKNgMcBs548VqXIdBUc4QMzr1++FrvOwgwUnUFJhoHNzONo+wEin3sJvplXJcm1ZW6
0EJeIaS9PUxcEPnpozsBlXKCAqH7Ddvd2QXIQlcedUdKbXdUnfs7cFv4X69OcadhJ+YZw87Cdhvo
OFVD5F/uXaRlvDwR7/W/Htl6yMmSKMdyWNPlQ8Hl5fqusjLZxxTSX4ttGNVq6Yk88ktOphkVNx38
LyOTdhtdl69i50Cq93SU5Wy3NUp+vqh7A7LwJhy/XHrLp//7ORccMy8VSqrQakBfVe1PGg20gxDN
bb9GtedF8Y+ZYrJ1AJ+woP9Kblg/7HyC1Vk+DI3njytEdtlbxwOiRxTcCWRv4FOt420XivwozM1s
JMpEKtMo99zs14aRgIKP8aGYt/2YGX/HsFH/kKdqRb8waFdlntKiAtN8B9i6iWAIBZ2tb4S8/0LP
xnCXJiJHsgqmRQO049SmkkoJ7DUyYoS2+haTiMLBnE8Cv+BsPRpImOsPCL4JGAjZ+NyybWAWL4Ss
HfvrmJhH0D9Oc/KiPdBU+eaEb99mkPdOk6e7Tt+zgA60lk47KSPGyhAPtPK0cbTBSu1vfTXr4fjx
wv2jvbp+AxiOgOjshbTPWg9zxirt/hcmT15Ukc1G0djh+M/KJ1k2SBHpcEUIEJWhB5Csk0PytS8g
B5R7Ms6ELBWjS7L+VkmxGpBDfmDAP/nH+M2QGvwIirPDYTBu/qe2e4zxqcZBueaVBum3ABOFuLi6
TPO+gYfaPsSNHHNHCtJ9ayhutWlLffzXCGR/h40hCNsiRF5vaHecjk2o1/BX3WTpExKVTGjaLW4h
mNJXWg/2oPwfwkgTzIq1JV8+3ca9hxs8hXYfB3aEzrYRFkA/K6NIoV7VWwyI7NRr/wVL3qiSxIHx
XkW649NbrV3rJhPMP5KCvD/4E0PesgFPTaptSTZj6LJIGQqXEUHDvGVk3XX5WiMK1vi6q561lRwI
6Fo6cKHJoHbqxjQqaxDfouGr+WWaWpecsnXfsK9fcO5dz9nkRUO8K6zBKzwiXxLXZTLzrndAy5Vy
W1Ty2+pG0JBZg+JilIN8TCPuarRcZF64C7McZzsggjQsWyHla2P5UGMOnOHMV1daf4OOKksOtdsr
EX2bIECUSPhnyqObsNZ0JXuaG9skvnXhRhBM9L2nOECcMqnjEMvQiH1cqjxFd37J0WeJwQ0/T0vo
Sn3ffTZdOJBIOFjnrl7vAgqJxdvkxz2ryy8q2QxSqTLiUjz61GcVQG/XQJqMgLZgVgmlb1lcZaWt
Do4Nleo0Pv/ve+xZY/2qeJQLa1vhVL7nfYIdq2K3zlBOUlPnUgwgITdNVcDLPTgxU6fg8wmPfZyg
JxCJSvap9Me2Av7CzvJQaV2/u+2Vfoeirz6Lc2ECsHv3/r3kwYkAQn9GnBqqrZS49C37jV6n+yUR
szKgrv2gJns6sZfQqAm8qmNW8VHpUFoVnd3ReVNISiPVFnE7XEO1t/md3P83SoWWVLqUO8Gdba7F
yIMrmHxo8iJEu+M6drI94/sZhZ7yc35z/9s9YRqla9yVSlWJvTrWefU79TuqRdTtKGq3vNcg+fpi
dLgYG3lUxli4O1t4p/C79r/VsV5Aq4YbiBw7ROqa2UzsHawlHmtFIOaEFK0a2oo5AYC9/uTzc65d
P0n4t8J6WFxfZ1t+MIvCKVYV5Z7EGGlV+HdFzwXQAES0oA2yaWm2n6pERY88XFleul2p0lsnR06k
lgxKfWBoQzXSenGfUkxE3Fb0a+WWv6HOun547v8wtFeYxaO8oB+hqEPggs+2Lam1/PzfYRa35ZEo
MzlsXRGadE4kjVnRRfZ/3DQvCjPCmGMC3aFN9zvBmDIR9Iq0n7rmxyz9MtqNc1mkLeuDt+iqKB37
/ObR0ixLxNiwJ6cpl1wMMCWuk/6eWtAXcod4v1xwkCEmgPnZmfnFoJ4abOPOc6h/wu9zCY2g+hWC
+/FxmoCkiMDGt6anzAQe1dJKWKP2L0V/6UtYnQGJe1zMJ2o6uRoaJKYIx/on7ix5+E4T1LFLhUzI
auBJKeD90qMOQHKE2QNZKtyxJ0W8q1xD3m97B98jln1kZT8OHJFNBevleXTOUwwsq7lOSoRh7mf+
WpfzuB7hyyoZc9ZliXPdzGXLXRAwDLyV4z/aDdcGbQX7Uyyu2rYt9Se3pF+jLULFMK9nFsEvt6t/
8Q37QL8xTwlsftnOlqcwBu2qDTc7rFoAGVmN0rBtpux9ugYAcrInOj2QzNlwPJH+v2VEowRNiNEd
wky/E2YI/jldfz29o3SUQwJypZUHLoV3ZAyaETPC/Q9ZO+xPnvRrS7TvyD5a3b/Ryx0n4A7uTJxH
WVUbTHJ/c780I4YmbIwCytr6wnsK3iTfk3Jm95t1tFtbDPqNVZWyITpEQZ4TnUdAIeiGWmK5NKCI
elMY+6ZwJMm8ujI5qZf0Jkw4gzTNy3/BAbPU25/5jZ8uyyidA7J57WPOTeIijUhvwwaZawetnN7A
2X9MpUMxjL3TJ8/L1etbgg5IHCJvcXbCQHqHw+0Xin3IckI1PiTCPTlVVyc05YvsluELKs9AjVT9
B/c7FEk7HxO0CLapHekdfPiRS2IKMeDYYeJgxgM4RhM4K06CDdSBNjxiRPv/JPHxHru79s/ewDq9
nZQEHRW09ucBBhDQoxaoIDz4MdA2uj6ZZFgrwz8wYqwu2WGwT2EK2T56/zAqeTu7k7o3vTBLp7hN
T8BXtv6rEg0RJkumLARyV3pEqw9a4brIjWK+c1fxEvMpi0BGqFRftH3uyi8mwPXIw8AgRT3f9fc/
5TuBltqtzYHV9PAabVXj4qdptrDJopiZhrdEHbyogdzwDAuPwhMSuwcUtS7kfddojYfdV5ilSPWz
qTuz86nojyQkmLmKyi+LTJpD6+QIwKlUYgv/srfEmBcUSvUavXF8l+Q98ttAgVnq6kzi470EtV0/
oK8ibVmebYdlQlxxyDYIKSZ4jKHie7n4NApP4cJoYR7nuDd0dA2wfry98sFeiZT+j4YDkmUzHA+T
aze46juegj7BBNNiGDvSwfu6SNeY5Ob+ppOkRO0QKKi/GeZgfMh6r0P3/GQ+j2ahB4aQDp7Sy4vB
kIqCPDKGsqvh2jiBWSqKOKLZRsxC1pcD5tZh/HuGYlYge31drdsya7Xc4wyFjMJ4qApLRWTBZk9/
5+IHuRNs6MEhoeF0ZWzOlpf+yKIVhWWwmNsxnf8e9qg7KGfFyVC1Yo51s27JtIYxmU6esF/+XoGh
5LPyODmz/ApawxFYrOvS3bH0WwqMTF5IcHsMIAXrglOJ8K4FNAp8jHCnAlKjIyRW5P1VJHeSbMm2
Eid2e+0hUUtqORely7aHl14nYNYazfapqh9DSko4djLlya3EVS1pTitN2ygXxkC5mNiTmc/PEjuL
x1GS0bAP9ZkAuA9FTxuI80JKRkrpPo6LUvWrWjpzGw1Xud6zwAAaOMCW+k1Dl5k0YyxS2oAz1Ugu
VvIZ6O4TFjZIfdfohf5hw9MJxW4KY+Aj2l3qW+di5fwt9hq7fD/Pa6JJSn5oFwvnbs4s6gj0QXy8
Dth/Paot2XdzpVOjzMr1GJm/5TrxV3rya9Kxo44maVDVb89rWroH5icDuCqcuJ8at5jSLWag1PJi
FLo0hdnPwjFcqvx59k7HyGYCq6rP4wNs968BYWHiTzUv3N6nj1/lqlHOgIIafjKa1D0EQB7RwJod
68FdC4uV4JjFADdAhnB8H3kHSK154iTNEkwXFYgsItQNaZQU6RVq7+FNFG3EabI2lFHuCp0Wb2F6
49kDnujL6nW/cwtP+m/MZJ1Q2NtMJW4FAMBjRuiRkvxlgp+JIlu52bySqjyFbXNeUP8XeU2FO7j6
Tsb5pQmGU4JZkt3NdIghmSyRXfoh2rvKjXRReoUIKCfVAHf/VS5kGfmbQ2q/5pTyj5nnFNk3mOyt
uxDQlaNMNFMg4cKHCt0xshSqdYTnCmTuWudFNPkvELaOLwpGuEnxsUJut6cMCAjaUMnRkSHwoYRu
xNofcmeI0VzjV9OqYhc420UNwGc1El5iLjn5F8BqFgv3PsTAxgTOvE7xCY+sRsrya5ZKO1g7jj1y
yB/gfbn8oUMIxspdwyA/aWORy86DFCOa0H+MjGSzIcCfppayqKk2rwzkeLuH1yRV4mj+wE/9vPRJ
xj6p9JDSDUFfovO/SQ1NFODUUO+jnWVnVuqWKSqeL3EZM4udYzR0bqS8Jisw2+Hk3n9MYgJIPV5k
Uxvo8GjbY1qjXxhDkrI7avmZtrFTdDFwkxHyGtOMPdDpRLaQwCC4teKOtD92qjjd1dFZeYj4xCW2
NmtTqA1xyPqyvV3Y+j7FLLqXztdxTb5Vmf95DSSPgLA8dDwCoKXXz2PdO4FLGWDwilKD27n99I4k
irl8FhRyTmho0EzBX1Fh1QiIutY18zrC6msVNTSJpzaGVHJO+tyhAXRONei5V7dv1fuqpgpH9tqm
9JXUDTc/xYiZB+FIVI1fTnA3m/FpB2jvruhbxOn6dtrT5hoUE3Mh/udqvEXXJxH3uXqfBhodkYk5
z4Wj1sVPq0g9PfF/7GQwgpE+5GoYmY8vvumDYtRHa//vQVl/bUK/Gs7nJcLpC/7OMJfP1SRiYvFa
cAE+8USDC3Jdh6r9A49EDA6lkne3iXyRQc/20QcNydZ5v8K30KtG7fA9HEN2ToPzJzWtocDDuRMT
hCz71DOFIalc2yotoL8lQJgaa7UXDpluZh/UrKIN/lvIz8mXtPXaNyTBaMGpq34un5SZ00kawU7w
jOz72ZSOTa2Z30dBvreh2gCDhN4Nw84JDse4yqm0QTl3mSvXe3LoEuZ40wt9ZjxweeeAWG20guix
RBs2rMSZYZhqX7aKHGHH3B321Io58MfgswJkf9m/zMxAcgEgUDlrHmoGzjHyNW7kbjeedKJEsX7U
2p8dWnAddaSHkFEA+sbtlceE4ijwuMTvntBmyVCgBHZ9Ncz4QqDIzxoCFZTvo3csjuOF8rxIl52H
16m5+PaOTuRVcPRp58hynUajhUzdQxfv/BYnCS1zKHQDrkt+fIiiyJWYj+XDQVos7nOULEctJ3f5
2wfi7f07LXEgdkD49WFBvWf89zeLNagSZWnMVmE3gw31TLygtfU0H9DcASvF9P4r/DGQKeZSVLgx
009gxvrTjP/qXrUoyIoSxinuILZUWriViHPsDZ+9CHMlmii9PsUWh/x6+JRVvUCJhzjE7L6dV5uK
O4Ja7eExoQ6OY/V2eeNxhbFVKySmO4U6C9etcBmnqDU4/YiJ/zRarZDW95635tmJf7ExwdN6X19q
wZc372ijQp3BVzEtym0m/hDBa/3qc1qnn8CEGeyrUvnBFf5K1KhzO3a2KG1Mb4fRpLg5AhueUFPe
oHaqQRs1IQ3PC9GybS+xadU8/wJc1aY9YQ8ISiGC2G+5p2MYBPAHmutRhmET4/lUHYJ3AMnm8jQO
kDUJRrYdl/vzn4n0wE47N8KxRelJtX/+9F5EftaNkT6SR0jd8CsfzXXB/Aj2MJ5XII4ByQ62FEs6
VyNQP0Oc96KYAg+msLnQBmBKdK7yUdpaNkb+750tOQIxoHWLI/0hdT5zs66y7sYdwNF3I588c4Sg
0Jdxm//K/9ZpKrHhGkbXHkS/Vf0A0WW62FlPIFhMzF7ocCk0MqvM7kGnOhgNAXOYpmFz/a9e5iFu
bdbl6kRQ5Y/RocKUcXyjZs/gu7BBSsqrA+QJlWa23fghYx4smi/kkuVNEKDDVkykVR7OHgM7fAwH
Tz9JgT7H2BanK3YTe2Mea4zx+Z14JdXLNomDYvNGc3as0Nrl3qbqgvbAQXjDu8xTI4EOQUq1Cm1o
zXjzIDmHiHaqa+LizZAFr4QPHElzez+rMrIIJ4GuJq2ZRvXcntsvtZ4+el6UkSQWwEPNLtg7hK/L
qs2JxZjxHldSil9WVgqpoKdM/rG76mZrre/mqWI9RUkmcl8B470snBaS2NI/+pi2JZWUmO7mWBdi
TeTMN19fd0MU0DIWGYzleO5HcfG7VhoO1/lI4OICuPTcAxN1ep+psbFZyuuOporrIoZe4QIGfw1F
A01U9ghcXOgYWukqBg2XZR6d+jmKrB2bpyV88Wp2UruB7jXoPKZ8SLZ2bEw/b7WQrg2S52WsiXf/
1aP1lLQbyWfpxYwu1zSIwI+tSKZfZaJsNxbRITObqBARe47uI1xkRpFahwwaReVj25hw5MBBg+Ho
sj36DNKStP3GlVyba01sIe3DVirUhxCbDlzxqE79W/wpZVoaCrG9O7NEZ0Udmf2Bln9xmfT21/vw
deZWV8NzM+NkbAqx1KzUV+zup0XP7WmZ6mqNQVZTM3+7v6jxv/ErzWVDUpKaRqhRfEg+dGyk85Rt
kxJSvVVJOYQP/1t8gvItycjMiv08b+04hrWJw+wZ65TR607NNdfNLjky36PQv+dmwf2w9qIT0xxB
PfayMmpp7mMjz0CathfAgbUcUpYIiK25DJwHvIAnPnyLctjnbFZ+bHtPqS6I1DKPpc/HBKoKub2O
eq7YifUKbZJ21klwpd+dOZEF/JdtkGE6AgD35wv5LJLXcUjuhf+pM/4cspHoS3yRg0qquUJNP7mX
oLKnbhQGNeMHdPwhRBM9nv9Tjv/ELtDkISyygYLsqLEQHM2j9dT2Xbv57svnvIewjvzAsh8ISaae
K4GfHoKnz+c7eHWMedgJd/Pq1J1Jc4D05O5JRowd25l/LW5yWb7dAaxKJcyc9o4Ui4Hr3SfRXfb9
WIpHzG2L+roS89RyoBOFlj1/k8utLq75vYinSe0C+Go8c1u5QbpmjWUeTEg9f0hgbA6DPMHtuO4y
QMmk0eqsn8rKcxHAfojR9ikoBwBYhCpVQ3OiXj+dyrOjFqE6JEjpXCUVZYRTs87U5i/oXFPnbqz1
3eN2KRIdNX/d4musfgqskvxEt4RIl05cl4qcLX4X78wpO8vBHeYKbTDu+fIORur2yOfosjGO4oqp
BelC/Y/M16dwoFfnxa+CMPnpdXFJ9+S6ChFG7qikR18F/GuE+WNAEG6KaB3qbh+LcPc04nNrtBtd
z8FGivdpeLDVW+zESae8ydqvQMd99jc+Mq+qo3WLtTcKffGWVAwIqVNszaebOGHVXGr80aY+dAuU
qXJ00z2y7e0mFqAIZeMToWU69HDAVlMGowE8MXr8fqsqTIFtw8jC2wSBLn+/laXMT//9/pcSI7ij
cLpd9BiqQN/tHsnsG3Uo3oY82ABXyK24Dcg1fLGL1qhi0Mb16ly1D84L4bfgjya+T5AC1BtVJB6o
EeGm5HpxJ9oKaeC69Gbfw3PxyylQhhp6NQFiJpjZUitDi3mz9id2lTbuSBX5HujQI11aMGwSy/9O
s9b7gmLSE+kV9oubInWDYqrEbF3uQnnQXMPJnp/060WYilFk7HdRQcL+EGN+IRr990QPb5LPWjhw
nV12sX556Q6esTtCY0/BdbSUpe/S4EvDZo8yoYm4vLJzWXP0XDh5gccQQB4b+tBuhf4rWq8EMBGl
G9mbyo3kqX4+yOYd+uPPAprsPB+br8+lPaToEUYoB8jUyuy9jl/P6fO4ACQt/DgW73DKCKHWbFj5
Qj4vo8rCnC1hms4d0gxRgDwabXS7yBRcjwoZJfXeDvbA1JDcYaPeYGpzn4ZfIvYxpyfW0NCiqsk1
M23gaPcoViNRumghfLfYA8/JTHYk0GIKZC53CxdBcch2boyMDCsVdjita55uFYUeitqAzimXsJla
xMGbVC0ncGmQpcMK38Tzz4+WD9lgniM7QQjK3NTz48VWQ/x9Zke5R1KNrjtRsufWd6LdrkHZkIF5
vJMyhNiH56cLLn9vw5RmiVsULuHWknnuB6oovLYzALtZiD0EMYubVfX0uy5UCpOq21D7qZdJTS0M
ilNSbiwKGUnF5eDvmOqp2PEv5XWDlPnNmyrKv/iZeg8j/XAJrogzeFJAwGeOjbjoGaHBCfzkBkkn
TXyYyZ2Ee1tISiFfdOKetMPqPAFSzQyRGw0vsb4HQh72F7lySh/6R9SE753iY98vH33rSxCN6n2E
pcrgfzBhH6FOq0YyBakyCRkMgwkw8YNuZ3rxO0pkA+dWi2yVw0ECnOvJo4+YGBayOpZf+KtPEs8r
sBF/oUEZM3WSjSnc1DfWRFdKjRG+sCWSpX8KHKLHPEowTZSa/v2jN+DTFIPSp7XHjjSoh+6y2IFB
U4pub6dNnHKMHWmvLK6rutxna0snAFk4mu5eXvhdq848/EXXyZT9ARWV91RQWuSRQyhXzkjoDNEZ
pSikyWL3tc9cgmUgRL4iZpXCflPoiGquHtCUe/vO2Qo0qdOG5bL+dVetP2t5Igyye7VfECEuFiAL
dW0gTZgLfHHVZDn2XTMUG1412Oxpem6NAYgh8H7Rjkqexom0BndBD17MNFUZTFkZD8I7SklYrKWq
p4WtYuWNMrNrPswucmwn4zdDqCQLjwhUYy20vp2Mp9yjkUtlvQqLxIBsqqXbg6A45WcI4/bCb3k0
2L/yz7U0TR7hnC1TGfjpg5nsDo/+FeLqD5mpPbzFltFFWF8Jv6Lfq4atBsovW2dbvl85iYjN0JXs
9RL7ZQP1MVoASYPqT/L5OLW2Xk7SMuhwhqT7c7El2y54T6naVE/wUrP1LYQK3469AM/CGNfrvKIo
FKxjpUBX3eC8bro2VJnr46Wu5c1kwImPWJsq1R2WmkdyxKcHxPS1jC/ok5JnRsO7f3hIj4/+/bMA
OHQRIz7+KHj3Lkg7xRIlntH8y9n+bDldg07cTJEGnBujKiAwv0IXNwyPx9HCPlUkp6NLxPVbwZ75
caM4yBlyzMTyR1+E2ROjGUflc9oaZdghGsqkB2PTM4/e7kLUMpThZ9PleB4p36Uu9feFzhX8yxDR
3ylonnUiBCFiO/lLUfJxuVoYEjNC0K6plOTcocC5MqPPjkMwqHPoe/F8Pg/1VEml4iT08Ihb2Lgw
ievTebdiFEJCl9W54rz99tDStWMHVClVtZlLbNLmfDYVL+iT5WRteMS47ERxxwWueeGbn0ced9wg
vOKtxxJ0CX0l3vwKmiN4B0sc701Js2vpWYwKRM7yjTuzfvr78ZxlJggMKjf0/Y8IPbkfzVa+AZKy
sVXbC/xKKT5Qm8Qs+J/qpjArC86HBp79ePLIyMv29aA3S0RlK6enCGRuDfrusTjqxGlj16c7SDnB
Ia0znQrO/O4QO5Er2GL9SmpgjOdt4gIFgbgPABTQkuxVPu50c/8DF/16u7M+rAd2rhhZnTkRwFf+
FMOE0SKODq+VBAxPfhITV1stYD5URs48DJO8B5UaGDOWYJlg7s56iwcGNcCe9dEgWGui0cJheMGz
iYAN+iAHsXIsajYU7PzrQtSeWEQA8NaPceTDM7Ywk2KOmRGeTojMB4KYYbUPrbyJnkcZLUICyyar
I/9+tpHDsec5Bgtj4k324jBqbHVMi26ClbSpWw5tU5kCL7/7wp6L4DacshltRljfTLPAp2v4fFgJ
sBT+z0onqbLFpsAlDVhm9obZ3x82RP+TUuSJFTPtf2vn0WX8+xUeDREnCWf1LUr2PBKy0JCDHPao
IBJ9ykoyxbyhRCjnbyiWoxyofV07p1A4kNjzROoLi64iBn9sj0rthBD3SxPqdnTKCgr/2F9sASNq
j0sO9UwHWSqx3iRjLZz8PO0FwHVXcYGolZU1OnzW1YGZqjwxRPm+VKqOhN7sqf9cmDsarF4M4Jnf
lq0QIHQmUvDnwr2YW5ZFVDxpwwUsSGOfoV3lwpye5ZSzX89CPufBKEDxyf6GItL3L3MXhb1JTTlD
U8sCXzwtT1YjRhQuT2UkiFxHNNeqVK8Ub6iJH5UGmBnW3fim7Nq58GBvEBmp92TUlw3wIJe4eNog
NDRndjmFI/Jv4geZwG15pfSEgo9+2+iwZU30QZLaUojMfq+5BEMJzItwycKfjyHUydfY7NPp8NeO
e/pDC5f2tYNQiWRW6KWmKwwtnQ239FHfrzquFKdx5gHOn8PwjEMXkY/q2y9Px0ujsfsHymEHPXNO
5bXH7P6x6AIIa1cxQKJy7pG1piOh2pR9wCtexQJk1HFutMDgsLd70GqmB0TQHk4v0BdgTbb9cx7B
9gNuIFMXDHlCbZ4PsYuwbqk4HBvnbJhuwSW61/kx+iIQxEjoMCctphw5nv8ZCg4luxJyn2fNuBFe
KrK929SMMJqMcOsEHGvbULCG/Qw7h0A4UHrlN/12GpycjRzd0+peQUkt3nWe2xZ02EVgluunsJ3u
RaSzrWOJPwo6Th9iMUIKg4RpblZmpJfxlr69YdwlDS+ySDHGfrPexUCqky5FgrSQoGigbxH23Gw8
3Xkf/sx2Cmn5lQoQJZW96XgvCe+VILdvyZbYx+p/xMrkj3BmnFrnN4T8FIM6WgLfdPUEv+x7dGVd
GQvfcSjWmpbZND3OljQQd4plmsLl3SawacJki3Z8OOcrhfJVkgH7gfKASmj7DnaY+ei+wHVc3EDy
aM5AidhHYilXvgI6iEj9LnnvOwRO6V+CpEFZDAAzGzMmjfixQhsISUTFUaFtfl98RDNbeoz9aoFh
Ub/E0l+PlZiIUbMNQYgdrlTb2jloDKckKGKBN0x55BFmuEMv+uS2qCU+XsVR7FfE13M/CEhrwO7M
eTMvBzAMlScO/aGT7bUZ63Zw6K5InK6wvCtbC33MdwGAh8ZQCVQNIbjYCRemJ6hf/BdrWm7vS3TE
cMMXINYUUgI6jP/mGGM3iEg/lmg7lIoSpO7U+ZdW+mCc4qWLIf0cLEK/rPQ4pX69OaPog+pOvOQw
h8uO4xkyIiJJiLB+5Y1djqWPa4qMfpNcIAJ4/vC6e+U0l77EOvcdWkeZPQ3zH90eE03I7sctnWG7
cEHa08oNWnxclA6AX/9TW1jxwx6hacKOqZmbdBKzFCWvXo+okTtXVrB9MPs2ExOEM/Yzmh138Pbz
8quVQIz9Fq62HGMkxReYp7IjHJTcKhOGHL742WrLq+eJOBiRf4FSr8z1tcEgEmfE8hbOD8J/9D5e
ITwN/Pp3WwHKHi7MhgQ1cWc4+j5bc0SE0z0JYBUiOIKl18ym6muzCACR/SUeemFDsVpwFdx0vmfK
goPidfXbEkTWaRYttlSpIqKTqGmS4JstSKFwrGc+Vr5texsZ/RQlmETZuEzsdwE+8yauj1W5S+uf
AXkjlABeKTt4J25NzTvebxZ65A+Ci0NYxJAS3+68hHtkT+PRK3qADv4k8Dr180EN45iTwkd/Y+5W
xyFsQMK2UMmTeGdTOwwcRQn5eMKMEsOsErCSALniO9M6cUd0hs4PcbS/bsHlgx6Ll6X2FccbgIhh
38Pqe+1cirNyKkypBVKyKjoYrqV1piiPaVRUSOIRolXzKWrozPyo6ruPFfeABcAFTYuIqzxWLEKw
xCewsoKhKSN9B60g36A/ZdYPzrI3bqRdKJhiJZ+IJWoK8hKPhRYo9t8sOD0ddySDsOJmCyLPDLm/
uJ988F3OVcExLZyq/x7kEa6MZte7W9JkHErpSV4FA0PkqFjzHSrd0SqspYzbYm3nvb9gWAnCBUPa
TumJuMHOQ93/Q8jISYGtu6Jsz4BcRCxgt0UcxW36MrPT6Py8MQLtXJDcLY7DsFapm8ozMAaI6Z9s
r9NK6Yg30MdB24kBaHu/U81WCBWdWbAsA44d/CB7RYxy/im/VtI3e5ywwxTkZYCap+nNly2J+Sdk
p+c/k6pX/+bqPnkh0i7s+omd09HTDmdatrZxKLz7oTwFA+NdEo9NBGR/eAE4o8lgR6YoTz+SycO8
qRn5iOw0tm/5jFyt9O6fh4x1vf5rd+po2YhogweiXez2gKCObJbHBPquclZVHJ/2W1fsdTZ1/jE6
gglh71/rqluzFmsI0vOHn3QNF4jKuUliAlSpubEDTCHg/hcJ0FsXdseMzZFE/+x560BIF+Xmdq0w
fol4BPA3BktGtfXVOK9hEzzFmkD0PV5S+EWtjJ3QiT8F9045bhdtuA0aFtaaBJ7FFOwot7m0Nj6Q
kaKJQTVbuXMYJ8iJJN2ReUAmx9iYJJbns3atWxL6bIqSWPEV6CI7gCeBFbKPNqBEjjrASd44EIID
+8MRnoDi/uTpWM8qXLrcwqd49NAJyFnFRm4LqnV2MTps3Arv1Y4tvJ/NwvjVsCepp3OvPcRpfx6F
O04nc9S8i2OWCZbrWW5nXqKDbY//SMDlvhmjcLask10kgEuvk3gDWOTxpMAlHmIiM6DkaDbDYm+m
bC8J50jTD/o+t08Dyvq+ex8lWn2eKnz6QdoVIbHf5hTJuqvt+fpN9heIZv9E7A3Tf3RowgJkKWcp
11BItTuqFha5AF2FZR1DEog38oW7P/fNw2nIaq/A4TrbE3u3OKMVIrEebuUh3sQL5iw5I4pOisoH
8AymDeckecfCQm5JCAJ6Xxf5cgjQqD7AJoVGYxKqt/BTXM3GD6CmioHeBVb4LRbJAJ013lkvHdnm
5qkWTwAXqA5AUNZVP/Y0O9FSKvmeAGPRg1SWHVoh3ogiiFXJLeurYfNsGBWH210cazmNfoRhgZIC
oiNdmpOlLzBccpbufbYzYqB14RuQLMbGvFk4h99MYbbKlQntmv1PrWGAqN81RSJNoVB2Kc8NpVVm
21VcUQ0JDTJvouhCCnvhX71xzgJtDE4P6Nue8n4wID826i3kPSYJsYPRgEp1F/8Xb07DMQaaJ9Dx
vht+Fghv8uOncpHtC1W4EFolS95a3bx/axlpkLz2NmQerpDjQiLUd2LRRQKN4dtYHH44fLAEV2q1
SHCAxsp0PzlJx11siaVoOXOVhV7JVhAWXdw0tZxOshzC2u2ZlF1SOzLvKczgHz5aIcBOzhkaORbB
axEreoNw3TY34ejgoLGHt3Aghqcx0itgL/Fx4YgC8yC1Eh2mDLf/ItUxEBO8zP9eN7FFYi6eJXLl
pm9WCEeAKN/whhf9ci/5zIOXSNug/dxdOHnak0Vi2WV8sCanxuQElpOP/RsbxZUtKlRXaccF4KLR
WU1iui1pyt84FdhkV+6nYQkDmvqA6i2Ubim2HgN5jkwrMgNzcSL1BUYaq0JngzIcqAcGYmJLfpAA
YQ+bxUMJKXePQOl3LAzkX7asMPk7MoUPstCTjqbvhW1xNZ2Nj4Zzd5VHbon7tHkHRS8EPKrvPR4u
+4ZYk9szCF9EH8TSxUjSbwDYWoh+g8w7hduXsRIEjm21b57vuUlP3aNR8MhZoq00ABlezvmgX3Vn
oxIDQw7Xh6EMsuNpxNvMGxAN0utpj6JrN+2vcBonco/KAzpL1aqAgFzyF8UND+IgV8kG1Zf03YjZ
hmfiroOOBy20yRAzlYAQBZNRRahNBlnixcjCchPo9uJagzs7Bw8ycPZcLNZ1bL7vqQ2AFTezocUy
w/5Eb02JV7L83Shdl1jDfGScQMG58JWURbB5hD8NFqDwMy1Lg5SYqd1n2Q0Ammor7j3E67OxRW3E
B4EizwW2ChTjXX54J18lXm7UUJDYnhsjyCStbUANnkR6bgvfOdtSltIOGmzGrz5ER+od/5eGoFGz
LpcdcO9VQ2VvNSopeaDETbL6TketmmoSradNiclHfuBYfCnZOc07678XDkzGPdpQfHVOy+RmPJcd
mIOi64Nq+NvYEVEk8XJxuW+1/wPOfVmCcreTgPTV2ok/7lrJOnH6Ripyma/67OXuu+uvUT5MxmYZ
BYDhukZETQOI82B1qLV2+jSFh7ao1X7sBCK4mme/rSi01yJy4SX7IvKdbGaYdfGFXTRYoZYhquHz
oniDqPMYXXt6nayW3RMTr3J3ZrhnSfbaSfXFi3WX2/pvaVCeJjJc5PVvVQBqp/sVQm9CgbS22mtc
aAJyNxwic5qBsnRgJ/38AIrUFAxXyuEfkDj+q5wFvejWnmJGr5iAU75U7Q8rUPj3w494ozP+lK3t
VRx1YWfl3/TPAVZg2l0j9uVQgk7nbQiOmkDX4BMVe4zzBLQ6VEVmGOIK072FcnlQF4B7I1mq/ReH
/MPrEA0dBZ8mE69lRA0upSqJ0jqFl5VfVSeAOPq/dcartGtGu58/PmqfoVufNtsVdxh3QEX63xaJ
VhQT33kB/3QWS5H0zOzjZeCkhnxnVkhgMDveH5sSWKl/Bjb1Gqg7ZZNCptxIThV/ggfWwLVcMndZ
ymL477tFj3Z0/osvM3s/S+XTWZzbVMoi4Rngq9+kVvkUk6CsSrukPKcL+aJa+GW0UTJ7j5tAAz2w
sBs6wSYq49OociIo5B9aqSsvsS3j5ep9pJJMsVmsErDZAhS75JgQiSOJQw0yiENiYcFhNOkbDWqf
4Q8oyj1Kofouo8eUscifc6uO1vqHHg99EK9BJ2SsM/pgQ9IldYzmtL0914A8nPkjeTlT/X0Dw0Ui
GCWD3XUHn3pahu6+614B6Ch5l9vuylcKLoUikYJ/qdAtEN4HY92f/El8GC/GnLCy565vAvVYMjKv
4UgAIjPHHN0ehKOTyNNJpH0PC5M4HEjjBBFBNtyTxkCRqfPjpSAJwpQGB23Z+HU2CqNhx+eYzqB+
fiNJv+DxbOhW0eKHSoF0kynUAHoJo6Wf8tDRgOFY6H1pXaHJL2/LihlfTkyIjn7OjjtV4E9fbISE
sJUNzVaSLBGzwnRBBBvEXHW0eH/ZbCaL3L4cc58yJoEuOMVTiZjc2TE4/CdX4M2m1zi32u8TcQ6y
DczLqjexbk+u44JgBV26QxGuArgJgAQRs47m8ATMzaHE+L4xCNhsaZ4SniXGgoHW3x1UXV3Pf0JS
nMo1hyGv/G90H+D4FpF9dkSQe9qz3woxH3aN2DeEhulg0bmebbowmHyxrj7UQzZlpFhwpFOF+9bR
7MVAZClrMLp19WBmOBVyk7HVoKmafYu+RaZDuAahgV6NUBixG6iUTx0Fy4AXzHdX+0BPN1SrES8e
6pfGqx0bJ8ZU44NoyYG02iOEmwYLUKAHXrv0MHFFhsgBfUsNA1/B/Q8dluyRGQjrq7V25CYapESu
2h1O6Ygub6qkCPFBlwLmablXoLaV2hxYeFM2WK5LljCwMtX2yZ64dCAChIZhmhRO9wne9PDdYbcX
eYGtHCUSYVaioWpjpM/PE/IlW6EiInkLPZhhIyAWf/1xYdN4YyaRi3zjt6Tf3iMa0DolY6YOZC2r
o2K5l5IM5GFv1I2PIHxNWKx549we0VRZrM5fvpt2Z4Ds41jyU8KwxggW2IkiD/yJWC3ITipIbnog
W9TX4VcxMu4xQ6h+yXFAo306mBTWqur9XD5sWk8OlFlKGpTNR4IPpQrDDeKsW6iZNpI5R8C1Fqfv
S5SxY58C9BnXI1Cs3JtyfmlaCiyAjjhhs4wa/e4dXZTo37npRvsT1OVPnbm7LHY9zQlMEcEhqcVl
fPJrzkdxSAxo2svqQMJdKCPwkBsBar+rfXSFC7KWHaTK7Eqb11Cq5Owbt9JtG03sRz/ROP8uyn3R
MU6MbLvoYbsKAc9S3Tlr0Y/nGWlh8OP/owU9Y/DAvDU/Rx/hyIn0dO66fuV440gcV/x1POdgo9s8
amVArmoJn9pUvgiVBFsgEPHOcJQLf7CBDzTpYj9Oza3mUdI3caI3JxX0BSApmf6hjhagIPD39uF+
52VoIFsTVhyFURfWQRDodBnhUsmf5Gi3tJss1VWUlIQQttt5hTyssnjuCLfsYa4SgZnmgSxHnQ2d
ZLg6x6dCnuzfNJ4nD8/dI5dEl6+d+rtDkKzJeGR9+HWBlxZxyRukVMTQW4aGnHh/1+TJ72WR3zaJ
/Huo8XIDI5p+2wLnkha2LywHIWa+qDe5016t3dgDRoJXprwJipE7n/m5zx5EBI1spMpe08kXGOS0
jJgVzka73SA0AlxPBZXoj0PL6TVhAW9vUXE60x+ezOzvOZxAZKpp9xYD9Nzm5+SpbSG28ntSNIY7
Wtmpb7KPImtLm8/oKJytjhe5PCUEAG6CpySIKula0RgmVKLJS8MGNctODhvkR2cW2sSyZK2Gccmm
d7SKAm9zEYfcOHT/rbNNwRswBRFQAKXEZa2KMAXWEC8oqBqhWOoz/i5+IAbeyIRovpWdk658Jeum
YRtvHl0lxbusfHYs3JFFNRoEgI1JLYQiuW8ZeoOJBOitqKvR9DjVxt9sb+OGBlMc9BJxuiA/0Gd/
qbl+1uPywkLMhPer6SARSppHjsLNZQDpmxqZQIaiHvaylZ7uuHh4l/W7xlqlKWdtItF5hRVONrGG
+0hf7DfdGqmBTYN1b6Zdl4ieIY0WwgYKVKOOgNxewhFyMu3gXIuP3Qemp0rmqYfVQwuiBXQEp2uk
RI0SBtwTC2Rq+6yUBEgjnOKqFD983QzDmXKZgv6KTK9BCHSGlxhC9O7KatqlcsKs7ePTiZE5nfYc
yBOxjFSu1lYuaHghjLmWnk1HTsghiwhGqSPbgou7G4ZXyXDcCLhtGjpBZgGVPIBxqirjGSgRWFL9
ywevcNwCuhgDIPqzgTbSGPNn5vC/FjTpWT/hBGv1HX7V0GbwIm7wKbE7NrEfptP3+2XEk77Zq7O1
FIYI8HZStEjp0TgpLgvSXwR63Z7OTl3WeNrSueZsMR3KEgmOfJCRFAURnExgVjV1tXJxRXtE+weQ
7uJBXpomctThNdan0F9sq8JYj8iFhb4uO9atjMz4UDMv7CveIxlGutPyWQp77gOtfaB6lsEvSIGl
koFeeukQcaQBkFidBgM11wt9J1Y5EkEeLcDWpiOfkekqkir5Jo+tlGFTugGBjWgJpPZthDejmpht
5lW60bsZR6PPHGUjtFkXDrCNojF/UEstXdPIgAN0mYqTiC0olcsDE8hBkB628DcagOxyQTWkQ9UE
IgD87oCibIF26vk52d6fJ4JjomSAI/57pxhxV6JG3v7eP7kl5mHlHmVnfsX9w2qzXsA2Cm1QDpQc
0fDy/lYwC7Wj7lDbxboIIrfBcFqg6DCku1nTrJbUWvHEmah2ZKyEDkkWBAnhyQOwUNoiy3yhvM8X
d+NKWcumsKG+8kMzY7sdomIXiy1JunQo2mYVVForFfWcrl50XJutFkjzpMBx91O6U5tk29z/cqy3
nQQtpSEHAk4kmxxrdGeZ+Dbm0EKEjsCNMykQEhBmU8u32gcET9K9lzbwFsNxuCFc9n7FYrgERuSA
BqU/1+Eq4eW/iGQpciPt55lOTUXEpbKoEmEOXbSMLkLhyFJik8XhbR9e88PMZQRyTvijiT2Jecpk
JVbbtiRpi2obN6WJ7RC2sC5AfmaL/uZaBnlZ6xP1pXvksMU4WQzzoDrZ5cMHD2TExxxwYFlKwGiG
5TekrB3sxVfB6LOpFW8NPMZ25txxSryTLsbNMuubJsH5tAk+lc4W7rLKkrARoUcOlzY3SzHKVdgS
uAc2rPj7PutBnzsdr/ca0zl7GYrcJhPHNQkDxWzB6A5WFpk1e443SD4KEg3BYf17uN/nCYCB2W09
RC5/SDPgyxj1relA/e//J8xXHJ5IgxZ01CRocORwXwCHeAmaH6AmADmbnRmMXH1yXXAa90ztvOmC
mNhKNl2Rg9XtSqP+K8Q/4rPS8KqhHUTFCLraWWUdQ9GNXeH5l67id5QUUozHAZuJIZjWZUzkjRYJ
oM8U2PhTIfmjSfKphb5s3t/EFKV//9Kf1JveEw1Odt+e7Pux1WZGtVaZUm3uc8ZCvTUq6xfcuBvN
/pru6x+W14CM+GaMewnv8wkbOsmUUBEIgN3gYCmeF7cFTtV/65h26Vc2MEh5LfkCCcy3qcXSA4oe
vOJ9CnGf+10K21GlogPny+RbxdvF7fVrNaCbHvFPyws1ozOxvPIzb2FWl3n3kdTMeSQamzkohri/
mhSpvIh9Obu7n0shH/yFzQAOTatRsfrdqgzq2eJieQHPO2rwtURK42+Jt4rwPa+30E1h05ZKau3z
hXr989Z5bEogYCApmJMG5m0H4+0AOZUCc5Nob1+1s3yNydSTwQghKKsVCRJjFJHXyEiKW4o6lVqP
lGGzX0L/bOhPp3RucK9gZQphmijWQ5b2y13dnCLcYNm7VoQmDSfWZle2Ob3cFGsuxnSUFrpOzQ/m
KxDOF5eSNBJDiT2Rup/67evKOFZBF1QWA3P6Z3XFL6os0IH8OcR1n/KYi7F2R6r72oiiYbAtXszr
ij+qVRS1heGOzfWnry8Oy8T0nWMRQUu5zxv1XC1fj9IlcUU/bJqh/pM+a90CuVVrIefj/LQII1Oe
URS0gjlJ8WdzLpwpk4SQogtVuvUyJazWFAbKlGeS1+ekpFbnJ0mGc1N+zPePVmo4B2V7tiXdyMmV
geY/U4UocFOUUpPbQ47PvyyXVBZwFvz6MQOC04hcHb/YhLXo+ApNXDGyUZbs/BrdKZ4gkHcl+dC6
VTIDTeF5QxHuzSF63Qe143AuTUA2XhjWmNdiaSKLNAsyq1Hq8ISwHQKtsu0BTyyFu7TSv7sYfmlT
DupoBubfsVRPD44Awv4homKUKRHL+ZnArkVAj4Dl93St1KMoqVcEaZqn8v0tGbCpMwn5+aoEDwU/
hT93mn4OF33RZCOGN4IkB/Vt7uAEOGkmTs93Or41agntw/x92pmkq4OSDgWZl0gBySgPbvaqypG1
0QFjRNuBW1og/D+LUevKhKxqTzgDUtpcT5h68SqQ0CP+nqrmpAc7RN3w5B4a/D2w6tGkhszlmLJW
oV8LcAKmOn1QHpZ74OBzbb4u9uxCFEDP4qKFMzw5UvaRMIB/czkPZSFSlOz6zYHE+MfZAcsNd8kr
iBsg0011JKt7SHXz6hCQTh+GN2cE9zAKUiGZwBRvQJX7tEbvMneF3+Zbbiwmu4zBgMQjWpmyUPx7
Ccu8lXTH8r1QgbsWXN5VUIVhEzVgBetoGIsse9YwzgN154JvLI7wf6bHWewlQMZmsbeTozgO6E8n
UXtT17VQZrlQfwOnKSKFXRRk5k2vul8CowXEuQHdh5Dmq5n7UCyWRV3ybbwA8+VX1C7zomjZ6A+K
I7yY4Dvw0OjTpHo3u7LZ612bQ4H8qqo98TLWL85pOV6wIXnpTvjfCyWpl50Hdyzfxy+jVVNSEgwP
8TR/LaWxvS89J9jZzbPNbFFayGgXbn57IJQ+ZI8E9ZGmXfv1ChWxay6n5dkgpUZ5xB2V39fUQhF/
jN2SuwzinaLyqSg3XJQtu39ibmkhhI+wf84xXGw5lBMDDlARcPxQEnz3BbTB9QF3Nuz+3stTtOxL
2L7P/2PX0nHw4IwSrNe4/gzA/si6L3EkWvXUYBr3dW7NmCUPauRqWUuuk4HYp3tNrnDAt6OCRe3B
XRW9r+yLebH+Um8opjgv6/y2niRchB/FxSCB/L35Q1a18jgvN9OydzlLTGGmJzZwO56ue4hHP2J2
LMHbwBSybMBqcjXJ1DN4D3FtHYppiap0PhTYPnw1G5ZrbqlBTL7yVHChkKW2efU2qkMOZw1fRxbx
C9753tni+yX0x0Z2FRQvloUyhMJkS7RGEfj5iscxn9dwrJ5a0WW0Hdxcbi46eK/oUF+8rILgmsx3
NmX0IhlpWGfEtFdjyaUwN5KLNQhc8bPusNgf8MsR151KV+2zAimMgt/seMCbSs2CPV5yai2J66PC
slbh7zNEnF1ZauTCVVr9z5fJt42U3kB4xJYpeznV7zARKDTIf4t3+M/GcD4ZftV43Z9fL668Gm2C
nBh+6QLQnCguyoLR6WI2rTcTlASTNR7G+qdvRR+rqzvwvYY3r87YZRBwdXEwMiTEYH56Lx/x8R7W
Qg4qUfx5CIAnYK1u9kIhZ4eQ86kcdGbZHIQOHZEKedaLf3tV9XnZVL2ZF4Ch02C8dfZcOQeZw9Fw
JRzTQCRlrH0mzw+IwFk5GSw81vH3xln1M0K74g/TEFDB9pE3EwN5SAzBLFwDr0mDJKiB/Gj4OuF5
wtQFr6xQ183HYnYrUm7EyGEShlkGUkIHt9Numx3PfL7R9gSM+m7qNWSw7IPOaY6Te98WsWvhdbsw
QEccrhFlkCfq7q9L5xkQp9LIrMl4ebVA30HzkZ5uzMz6DQLbSxpkkACXHQBUikM95FNUKVEBqtfM
BBiIsGX9cWkAr2r/O8ASk3l8Xh9s8Hxb6Rrvs+0mOR4H0wGPLK5QLf8/9qlK5tZiPDg8PGbufLCh
/1uCmbYwrow0rvzKAt4ddbN3QPgnQyDND4zYk3Td2WcZulYpIfYoJRO2xjn70XWzII+CmDeK2orv
/pbeByoN/+kBWMxAgYdnthANk+Ka8gMLuB/iL/W06Ef9vmf5SDLH92rLp+Zf1wb/m4atUbF3bzzR
AqLZHAmTNZaLNqwQJbSjkDy9PAxTdF4HV1pIv/hbbx2qgOsYsACOlQk0AZJfAi7+sKWbypQwG0Xq
P3qIMtRqbahm0y1/u0LagMcwdKySJoC+IGxn3pxi9SmDl8ppQUciMYcJxCtv6ceCP79Zx2JKTuje
BhybpusNkMmfXs7H7Q5m9VmZ1D37i0CvAYWQFhz9AFiFPzuaP2l278muJA1+Ur448MFzEpfeZ5hY
7PQIeW2JEiJJsq4eZ9Ryifea95yXBSXIBRyIexkcZagNB8ahlggn4TuIiesmRTL3jCxu9m76Cyta
L9RfaCDL+bQag2U0tJc1aRWGQHsA99WEEvJhWqxQKgagCL7tAVa3yv+fc2TiKCCcVgs04OtNA3ai
yFIP7+dXHoCLBtGs98LFjtz0NLoNvXCtC1qBLcFNXIo+ZyFcbj8LJmu6S+iNMaJ2XDCUUTzfbdzE
gvZxLW1hBZf7aMIPYkCL2GtQmFQ18BV6Kse58Y2JmmY5NmhE01TY4yTazp1E7AP3RYoH8+VuZmCL
UgRkSGITntS3TX/pIOELrc4IXAjdrOJKwHu/kmC+4O9b0zO+2JHGmNrYbosI+Js763xaIYoah1o8
A8Gm0XviUrIFahrbJngJodOYsM1G84x0xdxLQ1NnjKeYnzchX14dzhugwUt3JyToFaw4z1u2X50u
dD/mYuvGZHZGrg3hyXXNOueEvMkdNbiGUcmUzJvCxykRjWYSCLRQKU9AOcITaX5Wpla/Z3W2EmUJ
0Wo9rC30quq0vjI7kajv/RXc6Bt4jPM9BYjtBn1HtpePOqvW1voOIak5/+PTxR3KIzBCz6JSF7bl
Y3/8jEahnlzdx/OARKNXJuwVYtvwI6qN/YX+QYS7URHFiZDzUYcms8G9vyfNng1RBp06TG2ZxRk0
Jt404E1TYrWe5EahjUyRyltWZpmObGRZwq1k9TBRvbYIdNTYB1LPUoR4cA5g9fABhAUvICt2nFO9
+HmX79zr6TfQsoCxcSOscEehkIFH9J36f/b239ju7ZcSPFsj/Tj/Er4rmK4JX58D6ZyELjKhJRig
xO5BMEMjZtMxmK4wdMjOJi1LMqCTmv4Oj74PXsMoKSo50A6ueYnmSPD6HbU4oo01xC2t2UuNVlM+
WnFOdUA4/R6ImwEaI35d77AzJXSfOLQw8RuFx7WoJahK5cJWIvN8kNptxr+7Swqv6emiEDmYgEgx
93qOjxXXNvu13932qcUVjH4h4GZBdW5xochfoMwo8/6xZhBAiyy4WadX/3cKvJaicb/VYNkiDQrb
4F6JCnSx/pAdGsd8uq1pn988LSeK4Z/9fbr2AzFvQlQ+Accb0CfpvGNaNZpooKWxLFzyRP3CfFev
8CBa3ICZFlZghyEjIB58bOtAsDFBJ5r4Q6K6uGUfkILGZvpjtq3JuNAIX47tInuLOU3mGCSVbSsx
N4iYwOjILCaxRl2Ixyj6Vegr1HnGeJgMT77miVQzC5VPHr4RNQPFdqxgd1fC9D4Z4mKtt0wzXAwj
23YgOgW3gym9oZpYM5XasQIuD5LacwMdSVE+xDF5UxxW0MV2H6q1GjwMyQ5oNygl1JaGCvCJTR7L
9Vp8kq6xOo/vMlho19gxKQzJmHURSEOJVRWA3fn09Pdd5NWIghBTL8CdkbN/CdFIqiC9nS1f/+de
p/jn3HV1MvqHNXLk7RgGFB+vRrV8UbgDbJjO1EcAqTBctWq6QCQM5qKaQVZ2nyJ4fdSy0cZMAoiO
h7bsGoDMY3IYnzavn/8SrBBl/gW6iYBAQVSOhUhSB22qGDdm50oMRYjdAlhfJakI3P77T9s1AwLR
5sQo/AFUS2gZ1K7vukGStq4oizbT5a0IKpQJ8NjmAP9qXjvaJ92X6Q/AOBvy6gGvBrbWogiqg4mz
v12zpIsbxH0i/6BilCrEB1OYDqkBn4XKQ17YU++D6MMropvzHk1gjfk2BZeYeMBwimu3j3yYLf/s
nlBVxHxxhbAPTOcTRIc1h1ZcVDxHFwcdjW9ZZMxPnQ0ZvBYJIZ5ZSz5YUpdkFpNknskXyLAvKzZ4
7ZwU8y6jqL1VTfdFtG3Fwyq4ufe6STMrjQ/deWRh9en393ybeyGTdQBMTwUdLxXjjfcB2Lo2u2eE
bqnFL2jmTbRMh8txrgz2D//Cw75CcjQDUuObUixruXprf9lqah03c5kfarbFr5homPfn1WrlxOzw
zHzQGYI9tU5W1dNkRFAkDr62pAq0Gxc4LVpt6rlQKjIS/GDLK2pwXvjErK8kLg2JjUv9p7b5fx2u
5350ypJuyQ3nqcRaY/w3wGx/6135H8hK0V96Za4coGAwnG78ilK7/l0RaYF9HoF5EfM/MDRDW6o/
iSduLjkVP8jEYDPlkEKpVm08i3ZdxhmaG9S5/0v0kFwWg0EkBH0HFGj0+ZUiSuboJOorb6wCdBtV
GTj6FPnMVJ1X9zKwIHFGJS0QAjPde7mqmUtj3rpRvIbsBpQiLEEwQAX5/r2zhSDonKH+bMIiWuBy
t/Vb7+tQ9lITvPzSmbSNEEm+CHAb6YNjELQhU1wh59Ykm48lgedrRlHtXNDR1a9rnHoN6Bd6Fdew
3tJQJrGtam7XOeG8f1s7QGZaPxNbOGDsdjuwxs/Uld+AOuY+x4e6Ii41ChmB/PTv1Fkapsp5mwp5
Pe7BHpmd1YvDw6gxZ+tkzlvMNFBtmkR8a8gBhPXeCMA4VGgSeU2W0RguWwdAVBJY65zpSRILhECV
L7q/lrQTWUa8akel8U7kKvB0ZH/EbP6DYNufrMnGjomuhwRa2ABZsCvP3OqNGy8BXRgqW1DopUGS
i6gqK5jcByqZZpRDqpAJX2uCCt7ivXwHos0ctqefxuYRI9IZBVBC+damSeZOlFemXAaOa2/BxelT
2tMyPIun6XWEtvixHJ+vK5Q6+hpvvAph0czZUy2aK6IPiIqwftrXEjD1FeluBqCHx73ZnRc6SOaJ
+E+12/i5Fg1TFxuKHFBAp0fR0wVx+PoB0MToveFDYTFWz7bGtGwG2IUV6fqzw+xbDpMRC6tEdoNf
GLfxSBW4turSDHTusOAYWzt/aY4RkHBuez9IzbvYh3X3o56ll9MNWt34bmvP7O99WB91xCvt18px
dSEFcPXu+OG8nnq9I31pdIxysRcEnTNrLMFDPAi3P1tCrbMTnZovoBsv7/xgiZ0L5/85PRP1wInI
DlLoB/UTmNq6Oz5E7g5XLvUnF/Jx377ulWRpko9DDgAeGYXiHTyA3ZAZnaAJJWz1DDRuXYdiCPct
VIn9clGAhsTCGn9owQKaROS3IZisAXA6pHlWP1sFV8H8VjaYYQFZiSx4tDL/2V9fLGQHKNxJIBnJ
/eu6xDxcW6Vq6tQZ+R4KgQumtilImqLWtYYdQRlAvP0s5TGa/vMAiVDPc3lXj9tuQSKGD02nQcfd
OswgVWCTozAUbGB6xKiwxOkKSMdA+XpqnNGAEjClazPibE6tyRvtxx6GRrqE88ZTqC+317FLcGdN
nSTBWqLE8miZFpe6XX7O8yly+mWmM/6feOw/p5febVPKnZYyCC1RNAEvPKR5m9J+6eB8YzEGDxYW
ylv3+zMXEThTs9ie3vL3DhCPb+kaxT7DqbFQ3/XmJ0eDPV8+/aZ1nTi2LMmK1WRRjMlcB9kwSBtf
yMsHfmSGVHvftzdm7Wy2AgTYWPlDPAf/A2uYLdVdNbrF/jnujGNEs3HD/2YwV5rTf01Mb/YZ9oCv
RWa4fXDNIESAFOUnP2JCBaHHhGx2TeSUNYOFkK4cKlxFSYwEPsl7GUSfRldvUBJK/Qe3IABdhMvO
gtHmeKUvu9HDidRA00W18HBNty4XIcFDdotM+3QhM5uTSW6OF1SiR9opGac58xq/iArDYmMXUiDo
eTlsfS7Plb2FY0Lo4kMGQ6cBO5P9TN1CAfr6Gjx19l3fcIWWeO0AK/hJZ4l+X/CTjJ9HsiW5XvYe
xV4dZ6P6KwKfiJw0t9rsXWTm8JIOfs2ZV0dXz4YZVtzxrzN3ZoEsT2ShEi/mrSjUKntjbWHZEHUL
VVl/D7P6NC8vPFpUxNCqvahaWVCZEVsI20cCuHsDFsk3KKKoppqC35eh06O16/UxY6uB1V/IOEs9
sXYDokK8ZjvvwBmcXlXZ8Gi4/nro0ttSydRYB6wQpm+NIhGlXkaAjnlZg1QYwG7js9cbExNsCsWl
5pME5+OoT0PLXw7dtvQBxQ7AbWPaEvdN4BDvUnk/Ov2d3P1+yleHw3NVP8uLRLbj/DKnPCZEePjv
en5iU8sM8PMAwNtKTtCyCGKCmsxWgDV9tfSkWfIrBAOmomCw/1kt/dBclgbu4tI1FSD7B7AEdtYh
8S1fNBeJJXn8QvCjDycmpSIO8OHgloHeCtXZMpjS1e+Hw2GPViSKFkaPnqcKzwvG1iS0yh85H9ip
YI2BzQOJmLXOQ7BXItCHUEIz36rXINRXCOJzoY4K7CC9ZglWwdmJXk6v6dpQAsrCHXY58qCQLdpl
WO1qWyRDxHBOl4BRm+86zrEO/xdmXCuloRrFtp33deM767I0AYvddhHxjKF8fVk9QC6hOEGgHX1X
eyKQ2wtCpc0ddS1j88opRjt5s9RfpWdsM2DAyWL6M19ISSDfLf+kcXLnPYPEeRoxPArQB0g3mML7
9ZNCi9ostog/7A1mBhI+fHNVL4O6Bv0P4+BYXD8X/66lrvoFDAdHYOoOzlWaaL+wpihh8tLN7IpS
R1XCseOXvlmCT051lUvw6O8QCGGH0Y4hC3g9FAWK4koFOBJaMd3cB2rVv1QesLuuluuLpNvTnvi7
TgQVvDpwFuPU+jchhZ8KI3b5PAyvHocgO6HHAF7Mk91w8Q+B+i1Lv78LnbOxpYVu7z+65/mhT+RE
sWljBlNJVtA+I0KuL8j4sA7jbLxgifP0/7kZ0gYPcBXKf+xgH7ked/IlPSNG0gybc9H0c1J2MZ19
3jcpRze5qyv4w5Et+27gug2SmaSQe4704V27Su7Am9K6YproNTntlf/5jBGCqHqhwUkIOY7p7blZ
RF34/FGD94eqdjVEd0CX2N5kJTaR2FNyRfj2trZ7HX0jWHNlqvcKuEdulBv0oyzBkui10iclDPjC
nRBqVFzF0RFOIc6eJTWdXJe86E/KhtpKeHyeTVd5KbNl7WNgn2FqacJb3F8JEIHs1sdDbs0mYwtf
O9qNAn+QOcwt/EcJ492ZuIgkH3eET0bCkVts2lpkIymcVYndqBxVJ7yfMsp68H0YG/PjU79lEzBw
9PLg9PyQeWM1RZfFvvjJ6Tcx2XViWLi6WxmfsGzn7C1JRBaXn99i/oqI25XVE2QH6eriC+d9+HiT
3i8Uky1RAOJebtv1CO5UeYIxX9bUYwhCw7FDyjs3R8snthG4avMNzrTPN1A9dQk3hn0J9FjJjIkR
kdwhzvZ0LrMerK+MRVQGj88Z0f1hwR8AQiPjn7TbGKzgYBnxmkz8IkvlDqetCGBVqIL9ODnoFf4a
FuJo1TYCPubvwJZudZSwQkEBglj1NHPIPakoqBcSXDrOqLS960pB7NBUgv5xda1+d9USblnD1gvf
nGPMW0P4XwyNvT8hBEDp06B/tUF0L6pzldi2/2m6ibzlfI2JgaaUd1w+PUF9c1bp+gRfhrhcX3Ah
8meWhUxCWIaj+wM92eLF63YbXRtJb28Jrmh6SjvKGQyQjFQ4m3y4Y7UPDTfFUGQakKS2e//WVDeM
hwphjVR4+AwJ5IGZUyBaZE2xv0RVzW6it9551VoHLI5z5qdtzVlD9UDqDzhyFZQUfHHHDBhM2IaM
ZNb5CKYEGv4gSirwnvZUtZDIFjCzYIxELk1F/si1s4k+S61iKV0w7kMxCcUhIyN9sP34p77U7IlP
ZCwIGwAtGYmM3nCVN+8HH1kQQk9MqrMINiHN9v+D/2q2yi999kqPwwbuLy16qs4owGKTxv41Mmbs
mMs60b92NCl3aBw4QcLmJrVWKFK84kY9/mfxfxwKbbfQ7ECV10gn5Iip4WhoEHWE5yRIq7fMI2l3
xS0Hr/aRgMlZzQDGEb4YyDQsBlNYMIIXcGpu9Syo7PGo6CUbb92bFTCO/jfJliVLNrh97ATieMOQ
PeYNJ2YAwqZTvpczVt8Z40E5MAdhrAO03QRoUih8P2RJSZHEQkuZ0kJ6B+FtyxiTY6hEi8GiR4L5
A50Iuno9WgohR1txr05hTWq9dMqNFjJILeo0dSL8kGmpgEP0Rr73/ujCD3LA4bF/OBS7xgSqua/N
c+D3bi0w5oF0ncSWs1veZ4htuswQtc+JJy+2ybmX4nEjfJ6rpUbrnbKG7T7JKWLjsZAaWlBpyXJy
Hh9X20Dy3Id2SSjvES18iMXBULLz/BzMlEVrULf4S6+ymuaDHdkWOfCUYZKIBE+59FVnSkQpNLCn
TIe6KHGKZODJwqw4/4Q+qEe3+71ejwYYJESl+UcfzuSGaIRBfRIanPkw9YcDs70eEROKh/ysKC/S
ZDba7MDIw5799WCzMIl3vciengN3tPu0YSEe1vKMY/FsbXP+i5ngz6OzRp0pdYQvHMv+Gi/Z8L7V
6AE+LVs7Pb5IiRLKHtLcg39Dn7gwR1SWMhk1Xw/ThNfNKUI+EhJYGuCPOu35T6lm2PP2kaw38Phy
k4TlM29XSqD3XU2DjeMimY0kN8QMWm25A1AlGgfs9tl347iJxgusblNU4SNm4/Bfa1y/qMjMGz0Y
IaqTMc1+9ej8qaLbi/OmRFEf16gpqkpcERsBpuveJg7dctxXVMLRaD6fsSC/NcDKVSS7lxMz5vVA
vaOGXUrX9KlGRb/FIlhN44J7j5G3VndabqbV95yxl0EwlosYriSYWgZQS7gZjO+vstmO0ICfSVfS
uMkLcAksTStuai+c2T3W/5qZ0SbkqQmH6XV7zuQpqDHF7HVk98eKKjy+WaFF6pzC+GS2yvayJKzN
lozmFo7iCV0H2G/NE5/vJxe/R4bEPg2FOCtsxmdddzMMMnBiauMTrjQV8UvtbvINVnKb+FnmnT+O
5Lmtwgkxo1RTtlPcVnpEpulTtSn22S+yC115lWRiEGVtu77Hd6HdzCVbDigmeYAv0P6mgwIfqIRm
5V2khMG+5hMp09MpDVukb31BWVwvwATYgucXsjKioCd0mB288namuGeN14Z705meERvjWxO2PYDa
oUrDcT9x3SbFvv9iYQPIUcqjEyRLPjVH1w/pPgKKIVzN1iP3YtcVFY/TTaGzm+gfTo5D4WWQQl58
gi4BrFWAARpCtSN8X9WPYFhzBWXN2UKIXJc8/c4gIty+ha5jqzRBG2K94uwuh1FGj1tqwHhVM2rb
tjwTgcqPE47tkQArbolA8NUDi0KI2I3vtAO6iznEfIgqJ4dB6S+TytC0eRMWB6iUPKbt4/h1PpRL
x5CD8llsZXZ5onwioOrwx/7tHzV0thNOGatuJ81jR0jWWvCgn9D9XjeIvU4OzN1/eWpIR10ka/nK
vdj2naJtF1u39rlEzrO+MHHEUCx0MGZOUNf6+zzxo9VlFAFXf1ewMQFRubHlju5UxEZ39YuKHfAk
y04gzDwJ/MQ0b33wuNmUSGjHXmsyKentDio+1wVmYtoLoMERE+n6DaFPuizufXTu7dIDiArONdXy
8TunvQR9WkqXj3KVYQNG9oDky1JqpeYULLskKfntq/9ZC7PSBXMkCIKBRIIkBqPrA82CHW6HAWkI
Do6UVUd8jTNKQUmYPlVKBasHuxUeszW59CBhkay8fMVRYlGK6gpeZPuLDbn9+ybNYOiKeOp5nbxJ
QnBmQiuXyxFHIhiN0K4wq8Yci3u47T5wK2ly+DO9Qmq5osvbiOkCpQO0xQenhxTOc/DM5b1cj50y
5yCCh4NS/H9BU7S715UBbfySEiLlu1t+mTyQPBRh2bqbEwFRt+YP495dJYm1q8tMP7eLe3DUOVlX
6J8gZr8Ia5aiqKSYpb/3R5olQyYBpa7eWMtpm1n6fZ9MtxhvPk81E4uK2fy6nSPoPXI9+nHedoq6
8wOS2mXydCpVbi33zs6aEoLxTJ/PWIlKCkiYUZ70+WfNHVaIA0oPaojC23NRCFdSglKg+C3Hgn1D
+z5oYdz8RR76DYy87/D856WO6fVrRNoBeuGwbaPmewpQM1yD+GlWTY2S7z8gEuELKwhJdGQQc3Vu
B6GsNkAbg4tFmVsYXuJ6nGLDB1Dzg4OXc7AuArAviYf5hWyHQFwIjTwChQiXiLOnJGykjuNTp+ad
Eg3PoIgYyWwgdTsWVc2S3TtT0J8q2QaCrcvLowTvt5lImtUQnEW7mnxbKRU+o/3AJmzweFR7QKKV
MYnLDiJMzydXO78JIBGA89F+18PScq3QwvqnoF35daThjPQdgPheOxVwDF9X6tsQtIEkkeL8TrXb
03BB1fEr4kOJ+gyux1GbynyZlnqLeUsVcIo/35NZCP9POGJRFxSe9vvTz82QOn+O/4g2vGDssVh2
3eKWHNOrX5uamYPQV78XdjfAUjWq4PfVsA0OoJk1HRtNKu/DP+DkHkbr/KNzFcsB/SYaQjb2qs9n
7iTvphODQ/sGHtkqzQ9qMfLYDfLKvPQgwQazZo0sKcbnVyWVi5q0l1YRsgtzYP6ZC/0xjZZ8aP69
GEXCJ5k5MHNs1v9kAaRO0pTQhr4dv+tBfOG0BCgAryMJGAWXYTUUTXyLEXfhWMKEunpXl92Ha9ZQ
mmLeTpnbziz3xEUl2AAktjwcgBs+EuksQapw3iBP79/U42wOdbZ2DVV+U5L7BbzohvPOBsXgqd9h
PaRctbeH24lf1IYW5B/nxuYSCbP9yMXr32+Hp7pE7HyigDvWl+S6SXK174UMo4cbpyMsYRybvXzJ
MAcVDI5oSU+2mDhF+4fcLy3uujBsZ+IVqrX/W87QVKb5Sotxv5eGot69Aqdx7GHTP/KPtNB0joLr
AmkWcfvzcNHmNwKPSMusUY2Cn/nTL0Kyzyd77bRCGTvZBriyTIajt6KTj8MiMOMALEzK5gpXbpwk
DZuiLZJKDIWPH/vnVR/7NWPXmJ3/yZWb9PUwNz0ZlXq2q9HRavVzh53S2VPRlsKP6dW/aPWTGZ+p
/Xj5ZNRao6Wfyty+HUgzDyGTRsTgQAmHVoKdOcwkcYUNEWYXpuvB8cfPByHnkc41LBdvL6QJTCHd
JvGsHLTU3hu/MAvETEwwpyyfQwYwWM3uILIAK1x93ksDebDTpaWoi5t7Z9E6sPzfiAE5res35LCQ
/RLVDwg27dsDkE3ruy2vLtaz8xeVFpkXAqYeAmje/4lgMkuke+jGAZJjFR2gjgWYQFgJCYS0vL3m
SLD3b/818KUPJlWO+sLvnlxxmCvuhZqq9rV3XySsx5J2vGTd7cKpI859a2fNkqAFZSxcgZcoBY5K
CIU7fqAr41tF/HePGwIW9XPYc35jN7110aQ0z+ZqCHOYrjqjigpKREit5PP2E0Lo7XYZxMhWq0UK
nyLzaYrpOEenKxZlJXISyxNiehk68aU1RVfkaE1BUDE6RCWfxVTjX/7z0JzoWXrpcX8ka7dPkwUb
7T99nRSHkGDBFjiBkPqYVL8S3PEWYopfJlsS5LtPkAjqo4aDRC3Gak2bZaA3kYHsn1Cw0JMp6hjB
rPOfdv/27WAw4S7cAMYNSbDGAo0SWtH242JTkUAXEKyijLa5ssYYoXRKbnYJpYe5Z3cvDB74qBNM
xILaiezWYVS3GqpNdq/3IdseWLAh38pYUt2qtRWJGcEurCxw2GuTWR2WPf25Io5nlKyFQPkhFSYk
HE9bmcfI8hsgDVJ7MDluPzl12vMtlr+SP5ZF6BP4IarD2O7to5+3ZJI+jVSkCoRt+/yMrCcKKEeX
VaOsHRdx6iK3NiSWusSvkM5+3kvtc2qAcC56MQNd0ZgTJ4DugIF+6EXlRf9OWZ6emJUZUwXv2P4I
cmNRSGgeuHmm0Rr2LoDZa441d4L/3QYNAldnZr88S/2OhXgQ7E8lhe7NUV3XpLMTF+fddQWVuT9b
LCSkQUVgZMTVD5XhEnP8GSV6hDj/c2H/vMsCw7WvWTeibwQTuESnJGxzFGjhBwupNz4kynllb2vv
Ohw/EgxLL0jSB1NO9KFcXrwB5/qXIPAaMIStCSQ6wGTocrNwzH71GN2+NToBcyKzPEE/ZmFwj5AK
PkA8DyDf85KBxM7OGyCcZkcNCgkKiKQynIvBcIkax7Mx6X9sD4pBpg9WF8j4NwO6JD9eHwelSFcX
amrVWF8o92BudpVOaTbkxZF3yt29y0ZC/EgE7d6G+/usrrdADSresdj9a/bwGx0iJPMuzfeepfjq
90QyGLldCMg6eNfnw9XQu8AcjxQLtOVBd8QO3xOwMP2fQYR/bED4aswOsIsKBzco267VuzguqTS0
6ovu7Nanu7L53EqM+krD1BWssLj1mwDKeR8W5Ml+6JBhCHMgylgEMRE6UHjWmobk7vecgxWnfRiz
EHpomZ/IIfMgtkntwq4R1a1ImvHGInPwJnNX9ZMMenwk4Udh/vgl/qQ52361zAQAEq0xpZ93DrC/
0k+5cIJQbCv5HquK8nq+XJaDgP8M6bkUu1iW5STd94zqgtnhB6Tu83BYGeKTFnbXNBCv3niUtogb
eNIBrWubVanrqHr2OleO0zA2Ac93RPgh7twhVv577viy5ByXRRmy6KYRXqN9QNNkIqOCS/t4iNaD
6VU37QzEQ/mbQDmfjmdD4qiAq3I18RoPS8SZDq7ZJFEg5nnyiMa7yYvWOV587XQ1COgqtvSq1IqT
Srnhh10k5u8hWR5lirLLVI0tqqrsMTq88U5euVce2rRCglcwqnFpEEvsls5PsMdhutbGYPN9Oqwu
iwB0CAfuYdwLva/nWVD/HLerayllMYGmXgTf+IbLOrZS9c1c49KXJTfp9d0ozgkNeDjQQOfBOItO
xxX9ny9of0EF2tPxtENnyFhwf2ZQhTJv3Qlt+5Re+96SrP7N6xoVqT0NF8RnRN57WwjXPyO/Oegb
ZqPHbC1hBuhB1W5O4V8cEdxS3i0wyN2m5RjNFU519qVCSHeovyE7uZsYPIK5q/qIVBTT5k0DJFCJ
KVBuah4Uj29mAdPR4gPGC02p9b2ET8V4ypaRWwIYSKbaYiRuNubcnwlIQG3SuklWRiTUBr2ihBma
R+w/vddd/FIFJONntWvS6sTRk7qs6r2RvY7nuMxzPUboR6zp8ZeuC7ixif7BzSAA8I8bax+8Xl/C
xZZiBHpZNXG8cuSWNd64Ha7W7aC848Eybwvvgs1MZEPpD219bZPS5/RbS2Q9r74aCaco+Lkt1zrj
nSSQfUDPEnXZ/dklDCfmygYvqo+AIA5oMWThFD4H1LR27WviSydgsySeW5pb1ydhZS0K+HZbxBZQ
M0o/PXwRNhoDSCUWUGTmXoFfeBLhubuXizOhD+CCBSfnWrGtOCdsd2tA+0C31jJLA0WPk5QZgoTj
ihFnDAcoWLoUt/mNoD1Tfodi0+bGtwEw4gVgEI4b0Vsx8d+8O+8uJ2t4PdzGvnWAlR3PsuOyCjBk
AkVhgLWhJZYtLKfILRTLI5e9S344wVrdKIUHqwQ70tlh4wuW9hDEiQ4zsjetvoQSIpGlgvHxahYG
yeAeAkGYxLthUjBzHyGv4WZ/88eW+4/Ym+6SzkgZxqWU54ncI4Iywvd1gnoVdcqehkyzAB5RLUDl
rlkdmoZHWjWvtHDF7BXEQY3/1FEFAgox/Tn1lZSY9yx5ZwVsHb4e1yxGrq95n/ZtMHSsbH1d1+Md
nlY4Qe2pn7j0XhSjwAVOXhOXt1Xl+owZk5Y5Afq2VMgVGa/KjVjbtGAf0b3oOGgENCGzcEhc4qF3
KVZPSOWjFgXCFG4eXfkla/ClOb9h5HescEW1MeCl9arNs8zfKNP5hTD23kRtvQSf3MgwWLfTaMl3
dmH9Uuzgh4ChnecsYoHtwhz6NbudcKL17HE5ClLu9MpVhQvSJRBJ80MZ/VRJ2GTHlXqQsqfc+ErL
a2vqMI2Q6yQx5fW3BLT5ys86xiRcDDMgOSTx6/bE8INFLDuCPN3MHPZAGrX6QzPCLin4qlZv8mEj
6K6TDBSIYhM46OiMGjM50OuCG+AzqClGs6IVz7rg2WBYaFU+GsaSnvx4aV9Vph4vzES+6xFPhxlS
ScI9YP8598S6r9pxXpZ/7VdvtHcxVqjimzpt4GDE8xRzIqMPOz2l7o6NWqM73tpmMKKMyasAVJlb
SRY9Dn5ENVHNLaiy3Y3EjpwyGMRZ8sRffOdRhmuu5TXLRocyo1lAWv4gCb7R4COqpztM8ciN5+ID
sjBUdmA0cZY38fxUUypu5U2fnPaLCbuyidklpdtSWeD3BH38YeBLN0mhEPThjQjqPTs/K1+ybP2r
DXhIWChCopsBWuGfAbk1rA3JRXOJTKi+OOjwaIWiAI/teFV7117k9WVH6JfuaQT1m+XWwVPkjz2b
Zk/QbFsRNGMBx5mWtx4DJEFTa56GgirbZo3lzb+pcEk5RgCq5WUDRwFhcK98z0PLqtsGEBhrlgsJ
HsAa+xg/q7Zch3k8Gpd8kuT9Vpu51ptlkPItMXxY1DnvZm0b8RoZPuhQgMRpssffoI9hk7NyVOdJ
T7XBrRtKw4JLl4TVWXp+4Rhnsr34GYFoFl7eXAUDHMW6ysoRLbIPXaBHqKlrhC57vL/GJqmbDkoH
EzwL2SX4iNA3GkZVBhx2ZbcphkINgs7YcQIkuH+Pne9/i3Q2NtsRfoVub8rV7/ZnXVMDZpub9080
dROD7lxRGdwrDgR5zdpyP+5br6YOy9DTxsKFCc/sxGb8T+EvmiE/Ao7P8BXmqTdB43XUVXXPDoTf
RgjVqxm0IoeL+kl+WxQSaE4KDEgMAGF0D82m+5mNMbZ3KVnCSPJPwr9+6s9VSYGMazkB2vzfK8WL
HOimPQeNeYzYl4HZfy0dZGrgG49E+Z1yr4pU/FU0cVm36QrdY/rBwuahW+8WriHKlk4H4HL8dw4o
/x32El9J4aP91GhpDU2MbW5snS2EvcvbsM55IA7nmE/RBAxmfwCxDJZJ8Hv270iyidQboqNXRpdP
3d2IKoA9KreRVFG3GvMOZBsTMLWMs1ZwS/Hgk0I9R8HQaen66kKOa5ysuc8XdZP+WsRks2xtQa6u
AvxttmZbtpEo+wxxHPXKe/KpWUCFXV1VxFXgQ+6p91grQgJVTtXlndJ36RTTwTW8rLq1WlQ5ltpp
Yf0QAFpXeMInatzcevUcNNItnbVu4aUOjxQh+us1TSavybeb5gZmg/jSXUZjoXnXkFzYXCCreaCv
LBTgqA9bPmwagU5zYBm7wioCEwmSkPcfPCfJb+aJqzXgjzdVUzmcvhtoQsk5eFfk0m4JDQC+JRtZ
ABU5WtPIjNzE2QjBasWZeOHCePAujGRgTyzcFN8NdboybiW2Lbk4opLmXOKeLLKvYiOvik4yVJ3p
3v2XPvVoqNSOhN+WjJUCvc8EGc6sqkMKDrb9Z1LP12LvcUOqaqY6Xaj16WNRujhARuUBjHY+cs5u
IAAe/SrNG0b4pRjHYAUHT4Yke1TUsNOfUCMp9iR9JLABvDwOg90z8DqNHWUaCbuXKTtr8m2IyBu9
ynpgr5sPZyLpzmWG3Rw+ZPGGMybaa6/dm/T/uwx0Id5GI4vawgzgwvcBZzYFPlHVJrZmLh93YlYj
a1qXZb1Y9jEWfqKPHSmWmrXDgOkHnSXTOwudah9w20Fv+Y607nQstSOmV+c0tvwY8eleo8GwMypK
BaYlTPa2KTtSobqnYTTkKsf7PWxU29+JaQjugQZRjriJ+zUSG9XvRaqG2GvyYgFqaveYE9vTAIl0
QHeR3ke+gEpae2K9NJP2InpI/Y8cKK/etyJ7MT4Htt9MPfKqaLf/pnUj25IdS2zNCK4MHLQT2FhR
4dP7cCySegn0STX6U6uyL360Sx/sTearXDN3f1pRN+0+CLZpp90fZoRLiGvHSy1L+sghIlbQRujK
5nJJdh8CflGo/W5q36hBVyrRuSw9Z3lflqxpwRHBCPAqLQENK9GHUAUBNdY1KP+2HX3FKVXwq175
bHX/KBSecEfs0AyLOQHqjVBccClFw0pi7xyo7u3YCs18P7ErPvj4HxCLuA+edZxeZuT2AfGqsH5V
VGf2ZomcjpkNeyVHpB/S/spVNVVkSGaQRkZbeplgH24w/8eKJiQ5Hm3Z+lLDUHr6UGJqEkutcJwY
pgG+XxFEhl5ynVzvIDdqfN36F9Jz8EyFQccsHcntiVcsn9w2uJBrBmuBX0YvLLep/Fucp6CRpUbI
YnnlU9adZCA7zfyUrzU6c5L8CnPOm2Slx9zzgrjnXuSCRT0OCtulkGmDZu2LX59FN/6GzCyPa5aR
wjmrRm+ck61XrqLBs+oeIX7kudEPyFamLOX+2u2JjQiAbF3Qy13cpGoHUgcy3hq9t9+OwUszgJNi
BKQUAJzFwINZqoDrCrG7okiO49+fvxvw6m+iKyWNpivb2UdZ6EZBEhQzQsIjjVHuWTE3MBvNYyjP
n73w3svreBhNda57CL6on+S+O8x6brId4o5NBq23QMvLWyqWOi9UTAuTsA+XBqp0fYKRHYjPIxYe
cwVcmTTtPf8oY+GNt4bN7RXaQsv1rqFT3qOQquMfmzcZLNn/7cihh1x/mEJZXh8YNdZmHSgwIpsb
gmx37N5BzxRi9wF9IoVZJlAgMSsONSBHezLi+E6O2V/JR3T8lsUfJ5XM9f/EVc7LXh3sqxs1OUKZ
5DDlFXTzm+TOxGKrvNg1cS7Ni2N2ibKEp1zkaxLnKCaPO0VRf9bbcdYsw7ABA1sOHU9Cc7Ppap67
XM6R3BifhsJzv5O6BJJvUMBiAv8GPgaSa+duAJjHhddXqKZjuo4VSEGmvtY7YXuIJ14wSAGxURgJ
i5KXvxh5zTD7UXT0z29HfyT/CukT2LGNMFgbZZCGco2M5KcIwVjEJHKtQjHwbiouzE+DD/kgRLQZ
FlraKh9XPl3OgEj5vAybxxsufngTJGtTgzuHIBsbcaCIyOyP8xwzdAVv/p0Wsu5TrA5sI1CpYoEP
HwQDK4j0M36AvT0Bxzzu4N8u0I6YjV84d2yYvNRJlc1ggzI6BiZchjT+Yt5v9+eISLsJuKfEJrJd
yW256WPu9Qw3Ot7Ct7ZDdPgohPeXwe/fGt2+fr2Yu+eo9y2SPrtit/JqpRoeaRmF8DuTuQs0d41j
EIpEEZHODZQJXawNVqqXWhBegKZ3MW3qb8X/Aojl/CmYQL8pIN4UyYfXT2BLtVsLj3aENKqvTdMO
phzXJcE6aXEwSSP92ikIau123Slie/m0EEWYGZyI4kqaI/lMEgUYhRNsARvF2kBi4LOWqHXe3dEq
6irpK4sliQ96YCzzQOuZF2qtRalozQr7LZO7uCc+Omfib0y+pGtolX9MMrvTvRXwkvLv7OHzvpis
xtWZbiItl97BA70OdmaCDXBD0GF8tW2h1pjm+Fg13fzZ4SVqPGAFEQ7vAj/mUfvX+8N8NFlXolqC
5IctEOnh+uK0q0OU7RJ3t9yDgYemjzHwdXwWK/P0IH5JmudkjjGgwxvsNA97lRPee/oG7pdP+ypB
6sbaxC9D5Rao0iP6dV0vf089VEpy5y3BAyelLxJaUo/5CpdRPT2QNgz0jLv8vKeyz4VyX0IpFthx
S3HVVgm0dwjSig6bTkxZpv5zXfH51NftTnWue7UxcfEkYTpPUUPbrmwMWmYUNx7vpbrLkDXj+rcj
c38pbi8CYOJgA2vaf7IcVSb19eT8bgrgMO2TSF5WTVzW2zxFe1PvnRXSLYiZb9peeDXLkghP1597
/P/73yex9lDVVLb3KCtDeosk4DalERYgCH9+qECGIYAqKlmk9aBSVmRorUjFSw60fWCHoB9aJXSC
+dIIBcvmUAl1li6A3GZAd8qfC5SE/L6xB5ZCuBZhJlJBxb+5wjS+iTWlMJ/10xNyqDmvfVwMc5FR
QLRqxaJjzoAmcgsUSxk9FG6mVfcJya7N5iBCt5bA3coTvkwR/EXS3H6PCPqi4LShlZpPkGKjJh9M
ByjG5daPMpQFBGNb1SsP8loyxIxNyNoFrJXIrujVxHJaB09ii4/3dTQmlawIMHp5X4uxCTA2DZTQ
DSlzqhQ7D9QYb+yX1KCYUF/NN4d/hy3E6vjb0BbLDdsZQUHsDyy11cQHpffWo0m0YzyuYfEEShgJ
W+MQCTkkJfCDqokwZoEBF0l+UO2/Q6Mi/Qki0g8LZ2YjxWxpAEx0Fn6zRzpSBuf2b5b6lB9cjYiJ
ZX991U+sq2s2ssIR30ZI6uFIIXxBIC06fdSO8Rn0d0i9nppmf168cN20zNQA0uSsGD7W3ShmygVU
Kf+7p7fuQdmPOXb5cxFXDp8gQgo7JtbeypYy/OGFzBdDke6IQZYWiuT37tenxgBAMMxPiEfRlIaq
kzN1jhh/Mz3kQpGxPnC46/rUhhXbLI7d3YEhmFQiHVheFR4mYnR1r02cF+683KxXoprzwIlwYPKi
TU3uzmqMbYZcuLNiWGgcMio3QFobc5fpn3ggSg5n6uP5RzHNyFet8waXD3wb9EWWFfO0+SNKJzbV
GTKOeaT3UV6bWRnTxOJx2AJW32/Iz5HBl0OKz1KJHarB4LXH8iXh/GD9pmGs0x2d593X1LClzQtv
GRbTK7nDuUVJt6qEGULP3fepjk0RUt8gWs0nHPJEWfwM4Oz3+y2CKxuXykkJJozlnjtbVN5Vf7cf
+Dmh8r5rjY5rswyi3bTOR08e7VRqyppD27A/6DYL4HwJ0MseaKjt/DJ32xKqtWY9mq9qdhvb4nma
HCAjX/Sj56vPMu4j3HNAM8b1UDUH08MVLpI/wDZun97k7TFTYpIEXRN9jH7NU/RPoAsz5dDyBlu+
yOOJFCQABEw2E54SPjRUfc1BBLmhwSoXTPfOK0QiQ6MArcB0NYDnx8aPxdxQacnGPOKHfeTs2EdK
c/gx23TKHda83HFYzPJhui0BN5tYSlqkmI22xdk6Pm0KGxTDL0Qqo70mcZml1Q4hRHVykKp2sfCk
yCBym7gZPtfO/5A/bTJpPlwxXWSp6axWCyr7IgOWaxi9DrLFX2TumUhw5ERitvrr28NKEjQvx+mc
TcQFV6NkigHgBKJio9RqWd42ZuSf5m3eGELXFwVma+Zj1Co4wu/sWD+xjAAHeWzLESIfdndbsZcv
zK4eQrK5Z6iaIpPe+jJlX+DrJ92xQNC1wj5UJ83PWSzwSeDIy1sXpvIygSawMpEd4+V1HmWZqqVS
xJPkh0ZtDnFbom4HdpfHizsu6L/9ygKDlyJLg6alqQNZGaWNdqXUqqHXFXPlAGX7Tcz9IszjcbX+
m7Ly3vYeZGr6f7rS9DkDeIlQuFqPlnjJ7dVMWwQrnImhnL1W3L9PDDmXQ/ugqTEZT8U/xwsiwxeY
4fHPKVbvgyMFY86rroS7L50Q6+RSiIh3fLUUNazGYEhe3BOgfB/WwhBq7UOsTg/LH8rIVzoKFw4U
KAmhf7HsEwzXBfh7WYpfSWIyBAwfdhbKhc4TBNtdR5liFq71q4lSazCdhyrOcVNvY09ZqVsvgvaR
xgnaG5eCE8OYJSpZg2q6WwOdubdJXxk6OSbZKSOJdOwNMxZ+APpxuqPlHp2WfgjlWwtuxu0UOINF
0FIAtKYuzPjMiy3dUnV9r64nm4SxyV9V2NHNBI2sdfvXme5Y+iYyzVoKOewgeRfGJGKi2Vpa2ZPO
Meq0FrZL7y3NS9sbfEVnFReBEPCFO7V1QcEkWCQ5PjFAYjcabjx+HZXJZS8vnZBICYfaZEbHUoYz
RtcHmuH9oe/5oYV26zlDzuxUO9VRRRj/+I1tATzqkpiNGozvGrtP3HisUIOvoeZLJYpgBv/tFhaj
qnYkZRtSA28H0OU19OLnvhdcURO6Rp4ZkELmmeVgs7o3WxWJxN+iHS6dc+CKDEQn2fwlmCu7MnWD
MnTqJYtqicqWHoUmS+n61jaTOqA9RPkUmwNP/vWi9vJqdp1l4Hs70J+SJZzROsBlpj+NnemRHlHB
/2moov8wlonoqUC/l3itCW4vOAL/5nrhI3NSDgwzPgx6RdU0ZLdCvgfG/Ia/rMQdQaU6Bw1sXqpR
GdeSFPUshZwsu9+adgPhYCkhogoPW07woJ5wUVCg7awrqCWQsjNSoeyndQFVhdMQeRuUMVTfGl6X
ftVNHEocWl7G4w/IemAhjfmbs4WjFJQ+UHwHOvuLvQwOTSMTMZrmYY7iMPcrHZCXbAoAZ6wxfgUW
77//XAz66O8bJlRWNfphzMdkmX7jnQvxq2B6VdvfNQfMOAUEjZOOVhd7lOY4jNvlMVmxmFAlP2pD
l1l2AmpqaW7IerljviulmzdsrqQ4Oc5iHb0R4Sd3BLIYHcRfKhm9d0X03i7p19HPpqFwjiqJU41F
kRe42W1m4FTApGZ2Vby7s3ytwzkgCOpGab/HNLuq9SEMqSLuO7TvYrUI+VHPto5JQRXKrmDXbjgP
8MDn9ulGJkXrSHbUU2GrZ3lDzvspeUuDUms1ZHU9LL2Cx7j2aXp399YstUBD7zAtC78dUlivqMg8
kt0vQ5ZbUbY44+z0NfqQzM6BNpu6MUidMlyL0LGRQzUTK8ojlfDVf09ESFxo8IeX4PAwxvvRxaPJ
l4IJdW6ODD79brpmnodYoM6MwekAPkpNGaUDNDeUOe7SV8IQjDpbmkf7V9g4aFwlGfTDINUq/LtL
QUOKbOATBKECApWMpp7nb01c5ipcEn3B1VMHd6WlEOf8/y7mqBPxA6USTu4q+aw0H2wY88X2enrm
OBX2kmN67UkKM3KYK3YXarEMv320UkdHZ+JoDSLvmQssXtaRMbTSzg4R770Jh6lSYS8Vd/zQRy5q
sOXYyWGfzOmw7wad1PlhgCc2Uw3xTqekfWJjEvAjdkEZlK9ZgqEPqZtTIRUCcFbZi3mi/VCCWOvE
T/CHs+ndnQtl1EXZ8KIUAAe2ywGTscYrkQw6n5r5nlk0qOOY/gda/D5o2xnAW7Prb+rjx3SE5uLD
/5VQ/Z/DPKDd9Mdw8o/LtjPv3MxHVoXiIQiAJIWIfrY+z/A3M5sPRtQnCC7cSxouP7GEdBENtMIi
YRIs3N4w3SD1OCXWC/BzFSy/etkuTkaP+biMoAif+92LEStP3KgrfUrusEttP1tT7+rtMRuIRBq1
GuCO0bni0uBT5TWYdfOnFxoC07v/cwD5OpnWN6rfnyaby8w+dqM1RoQ6IJxh111e7YLDDGAsnIFm
bNoysZBGIY1O44Oj65pX5DV3YlAj59O8kimLL1aOP4X8Ul9cglrWm/JHT8vvB6SoOFlMVfLdjcrZ
MdOd4hRb+skZHnr5xj39XKfty0diVKGQN8KLEcmqDdDRLK8EzAYGHOcUGKV7m9WycRYBp6/aTzhl
9FtuEx2A3GDBiYGY3v28JTB/vVsJRcoBhjij9xcBWIDvzjCN9dQgq288TbWpAcc9s3s6O6uW195+
nVRJARJPese/mQmzKouUZRqIeZrkmghYOEKxrM4PGO+yHZiSEwSh5+nwUvO4Q1zAkQItH4z/Vttg
oMspnbzxvSBx69LanDolsoMuF+SHyK5w8QM9hnDrF+W2iF0N7VO3sZZ0uj2FA/mjQXgxLhx4zEcE
zkgYJ/58oTXV8hlQrpr/CoFsiJdzWIy2tmGOvXOOCTeQ8YOexeNGer4eWQMM3biY1sMvORJqwTcU
y2mB3CPlk5CXYaObt/UV68lzo3ARiCP+wIc7wXJ7Ri42cON1YYPBJvQRWzzrMcxstHkUMUoaddGd
QKzgKnIj+KudJOSkdnt+4TaT8LjYxyNEWDZAKPDBOhHj6chTDvT6Ix+Bl/tO3BEuts24IAn4S4FG
XwbiC9uQ4VOpcKtNjaGmMdQMeww2bpxZ/j87ZJGSjpIU2FrOsOpmifTGFmKtogC01mAAlezB1+l9
ZaSMS/fCiWostTK6hpJVJ4FqVRHK0OyPNZeGiJ7RK1qtQ36WW6vfy3eRnmWikp1RypZxV7EENARQ
y7vGMe4qhDefx+9084wHHKVUJ8B1UZ+YLo2cd0G/2mDz24XikKul0pOQ+2hh5Q1t87IjWptTlo+t
dKRANvhiATampwWPQ1QKEwlzDCQwYpRoeZrzVhRPSpEFaNgRkcfpVzhnhdzQGGAkN4vA34Ub7NES
7U8qIk0rhHIqf3xCefiprE+eSX+aOeqmRvo4TJik6huQf/+Fk8/GdKN5MifILcXHEmItPMbeIm5w
xgYxXUHPolihIXzET7G1FYJcNUjLUEYEegHFgmlzdjQGrdzzceuLKYITtu+9XC76NPiCJmGBAmiT
XI3dLHyKfPWIIpz/a2PLkDsL5dC912rjiPglL7gMf72KXD0ZM6ffVNS/zdP51bO+lIvxemsTtB+5
V0735TGREWkkXZ6xfLgY1PzRTQw+u9DUPcOTLoOQddm9xIRGPwcrsAS5Kulfn63TrIpPdFSTGHHV
j2kIHe6S+RcZbctf2ihsS8EeuFoHRmOPrAqPzzaO/2yNRzUSFQkjwjesa6jpzPbFWCbZh3tblC4d
Ds1BJ6rRjC1TadR8tFLB7AE6XX/T5xCGvXqmAG35poxcO8e7OyWpvJCSpK9YoIiHEFeyCTl1VhU5
b5HZfvq/QMKDSKMIf6nFGkSnEyoz0UnKHPJPr76ytvlgBDkzf9TVn0EwGojV7qoYquGw361by40I
rJEmPCBZPR0dOFU3s8YRaJusU7tLE5SpM03ZCK9m9esB4WYrH77yKzlc+aZxH5/4V16TNLb2qmg4
i9mgipLwNK5VCNxAFssXs0hWW2q1G3m+Zmb7r9vvO025mMJ4uq4iQlTfAAS/xod6HRy7PxF39E35
r5pBDixOQ0og7EYzsf26miBV8EVTwcygeTL8Hkp1QUtinDnl1aeZsfrJCywcqu3QqwdZ7T8gitvN
e8nu8WJawivY136BjNmr4uuSzcbvh874NSna+NIv66Nn3XqqUcnXkOTYfZR3UdfoDWK6LeULsqIp
qQwxczCdtpcCm0jJT15Z2LpSmIQQivPpdfp3zwCjE3dPMmEgrqNNXwJ1ililJUJA1ldFu+i9MbKH
7a/5rvBvdMs76mN1GFYVjpndSSA0BKIAZ0q5/WwaJZJCDYfPPoXQ3AsvV/rpG8Iq7jREpyxhq6L/
MDtEI3z6ACaw+i5dLOe/t7XaySO7wg3/3GZbknYr8lUCmujej49mpnr6BrazCRDUhZjTjshg87OL
2lrYR1nNUZ4sop5/qIWVEx2srbmMGjOz9CKErnU3YTAdpeWnZyKEPuKe25Y+wskwJaMG9Ftxh2ev
ismZkVdWIuGVZhAYHqGyKpHSCOE1qfye8GpL1g1yb4J7lySfym4RZeCT7qHmNc6buRZBgWHd1GXc
iafCJZzD80CP8r6gydcAk37JCWGKCH+0uBstPHizgI5rft+lKwluzfO6dVvciM8tRXoYEnDL3atQ
UUTwSq+uvp2yiN/JMViRfpjLZAdBRCmvWqTg4rxNyA5IAVxD5pZqp3EjWEsKdl8hpLxqhZzwlXcs
saqIPhp+0Kkl7z1nj6/kfTM+CIwslPY785FxwRIQPHU+OkGyY/Xn2tLUpwz+JOT3Ric800jvedk+
5TrvpBvCaOJCB4CFyl3VPg/VOvRpOJNr30rfd4eXa6QUKfvRa0FshcSjupgiB7s1I/pbcUamc7Mn
oUKn+7YvsSd4luQCSCR4P18s33mU+a2MvIiTTRT+mfPPw0vyhbf/+s07OLDcUVk79z8LSg9vjd68
PqdrByDvRB3DOU1loQj1g41j9LMNyurW877h6ib1pwZbxy9JNNEsFpBvnNnDtko1/ehfu7J+m1XR
KbjbGUVs8gKYgTWxUzwmrxlorVn3/0Pcxte83rkSaRavImRWmeSmVva5RCBrt6/5z7eL81zU1Z1s
gwldaQbKdd00FiidDcl3XJNNrdRibwoAPsCAGK/EI9XW/iaPZh+1oXpaNceQB79WIJcA/yOUFRn3
VmgcPziq6ObVj5SpS1bHsThuskrEY+LxahJ0Y66l2oTFjOxS8QA1QcCJyBTBU+ZlJ966Rzg0PBFG
6NTUEqq1MpnpbKhvefg+f6f9GQ1EOePKJsqTNZ2o9bQ44nHHVb5XeAqesF4MzKsE5PnmsrE+gBkU
TWS+9yBqOIIgPya0Q1/ravb0s5LnjQUcvD4Wh3n0xEUK8lkcNzw4g5JcagbPjlwSAsmPsU0++XUu
juU/SjDEQYQT59siZnSRUoXEz22yWK2uy7L870WoEk67ZyOZTjwysc5nRbGv8sREqkfN7kKv/QhO
mCEjiHM1MUw/X/VOVLArWJ/LgR9P4PaIxxEjFlXCLGDSTxfGTLBxyhFjgAVOwHffo1z85is4SsBB
1PYWEumjAfjgcucSmj/w6ZcZAQpLdJ0UhpD9onMc/ByGzzREf6zHJupIZcNiAU2EVvGCFaHuWh4a
44sL0SZ8QIOGVKizXfueSU+sywc5hbDicXx0fJPxqHD8LBEbMdSrE1m99IU3UbFqiGet/G72hZvx
vzxf+0Uzg5XaJvOHMG08IE3RD0GQXoR4QWk9jOhcE/Kczd7iJmClxIUocBnTP2kepzRob5j1UIPT
GF7dsGIRXrLJNrq0HvJUFzQJ0NmW9i1LTlodqlWAjM3gKK4wYel5FlhMLGi9kSS5NAQ1oCE1uSQl
DhUTm3C7Zy+g/q8+N5XS7AzJ2ZXB+IHkok4Tiu+VHy13CIg1mgQ28CZDyiyEZDdKjRz/VLeX/MBY
ACKe/pHC9RNsW8KOn16k2AqAmJbXPkUP4Tk808xDMgynFTw2I4bjSBvLZ4wcXUBnRO+dLUvq6g6c
yM0/BRH7Gl9hmr6OxuQkYH9yAewRb5l8ELOE8SMEh0XojXtX+k7QB/ROsf6MfI+EWBfO0XSjgaIv
rpJCoXRFzLxB+DNbtA8UzHafhvqzOPPKr5WRrequLG0woEfSGV/GGrgZmxg+73M0N+zFuGqJrSzn
dLuPRLdeEz9gNwrsSJpG1Dun26wmklMYdXfSImvvxpqAiqgeEqu3q5DJ4XFti3ZggCxItOLxnGVR
Dy/kBKUS8jOGl7FAJ2kiT13FrPIwJOxT2htihHdiO7rFV7Yno/pwE5jpa1LbAFjGZS1V8DWuyCe8
6ycxS6WQxwStXIcya1EDUqbyjXmg68DVo5HW2lF5OLgjjODwOFYdGzQ0UNefDPgQF/my1Ho0LJBF
mj/C5z+cDy1frNN3gDX8X2LmC7NYoWss3LtuaCgcZEaJRX1DygUgURMd+kjuYmzePPmE+WCnD5pX
Y4rdWnFaJ0WTQ9RPzCRPZtfz/9HCEChbhZn5+6l1ThmMiNtEzRfCxR1xsT9q4lQC/7sLtZdGN5eb
M6xQ2mHTetAYssdz3xdVZ6BGB/CEAk8ONR3J20Vhaj40gwmhtAsevvSZDMVNecxadyDbmVrNjzaL
YjAGnx69Y4Gc2/sU/0BunCM5LC7EuVbWBNxfBk+ia2yC3EGby8s3Lq4eG4mTWD6EAnSYF1GQElrW
9cMmIKihDf6RdAdGUrwytMrM1QiV7nB0CSrDfLUTBk3RpFTrcW8Q+6p1meKNT5fuVSmu6mjkz1Ix
kpm/VhSACXqkCAwu8Pgojsz/rSIc7QLcfahgpIoeTdGTmoqJpJFqLaIUy7DQkED9p3sK7O6iXOkP
9ngB22B+a3DeoNynAw8Nao0n3kR8xbsjQ/EuAuKEx6lzq+ipn0BHyMcvW3mJvGoVzxsNqVob1UJV
D5seld+D3eApC5nehE8aMlbep6KcpEU6/UyvbmXKvCmwmRBmBEQ3mxlC4Vby15HFW8/WH9oy71Fz
uHIfN+DdGPIc6SVhMu5X4Vehskzlct7Ouc8akCsw4wpD/zYrcU65kgC3G/HyeJHF9p8Fn/Kmic2u
gmbnDkF+or96+7FcC2SrDmF6rFOcwuQurAopX1WJP/YDMbvrTVHo/O4f/xkAWd1g4/JImRLYTgDD
ZbiclgHYTnByQl3dt4t6Ltg90EOO7fsEvNb66qMwBJnA9UbHD/MM0TRM3WJwp1ZGJY1vG+jFN5qW
niXyf8ZNN2pzYx9NaVKTmLiUOHYmy2Si5DmeM21z9ow3kuZheSLOILynzq+heI6CtI/vmWdlEoIp
dulAuOsWV8V3IT94XC93yAASITwSweZDOEwwYcjw2rOTjD6tDO7uruI7su7gA0zpyUDNlR3huZMb
UcLYf/xlabDXYXcc2rVYU5qkfR1jCpwUdwvyHzLdpi2SQY0Wy3qR5GXzrL7ST2YeDt8zqw9si4SJ
5N/8kxBvUFfZ2sjlbCJv1ihKtjAIF/abzwTnbm4zKkNW6fqzgJWyHeHOh6CTMVZMn2sjoNxNpa4l
QtYREi37Cc0ogkz28wzJZfqjDisu5XVi6thSK5QFG8Ab3Jxn/AhfzuuviHnDZc4nAABHzUxGm1DU
DRBAKwSmgpbbvME+zENs3AFszoypL6Jd+9AgDgJczg6rEfWgJjnCRvlUYNWTEmDcvzH+WpL+daLT
HvhwZF2NUqeQBD4TOAaAnl+TEXmx5AhFenMsM4p//EOgAzN0NfEF9usOH6nm0+SXKmy6vEA3Q1q3
vfZd4X/UggVGkcTlzfRZA2uh1cCBNPqR6KTDSSyD4dfeBDt9283CLwHa/h9iltQSKILniUYizFFt
wvWcc3FTgIc6p45F9kpWbqyk5Tie+bDDPirW0rouSSSrAKSwtmmWXYqM454FT6xYqGm4BGHop9nx
8KsnZt7BpM1QSxFgNdvptj3iK1hqlmD3nJlGvuNLeo7pKlMKvmsoiWx2TTrvmQEmhZaCxHDEtnAN
j2Ne5HQtZ1BpyeIqWAk3+EPTupvYPU4Yw69OwDeXYTO3CdSCA4hOEktE1Z5eBmbHSmzbJ4+Rnf3V
50F7/yepoxJ0laRmElolfwFlSVipGxYx+XyIv7UfWMQtEggQ6am/W+T6N0ouR9Uhv3qom5W2Xz2l
y8jLvpzTojbAxwxpIAjOTVBpFN218i9wqXUcYa2EI1wWv7RDYYA8/nsTsOiZegg5hdM6UPyqcejT
DyBSLkE/zz5XP1Qn6G9R62PmDai7y6T3g6TvH5l8Yq6fttfyM+j7sNyPawdvUkyk2IHhHKF8Xp+9
AvfJrEmlMzJXJVGkhhSoMAIsJBHg30ZktG06KFI2K95AETrKYX4cs4T4wlkDm9Jq3TwxkOa8YKZq
slMvDnzVPytqjPZExEdBQKHlBJqr2uM9fP+1J2IYy7Ndknb1gTZFGG9sdeen+3WiCCseHES9mYOT
pU8bKHjPh+6BBU3nQZdJpKX7y/3ukvdP0VWY8pPgsSWhBJd2BywibBDpQL9XLkaqpscEfAr0rQT7
PBr5YBnoA50Zyuvjqc4TL/UNDJIXzmH/UmyYcdVhs4XlBSAd6A/FsO2pBQt4d077GRhWW3ns/JVy
0tlSFS0PRw3WqgpyDvcgtGmejMycOS2J51nA3pgj7BeUp8nJM/rnD7S0Z9s6S3mG05XHDHrUbwD4
kiziNfhrL8+gogtj6/iruomimgqfUvtIJ3kZjIRGuEsSc87aVvBHV5RQ69X4RU0P45jE9suQkx3x
q7wjuwE2ZHexuwvWAax4OChQ14HYBnCiW8neyEQHonMQTIxc/x+7U6X0oLJJBWpTPwo/trHfTyok
4rWZi30dErVIMO27VxmAJaWM/SH+SgwPjd5ZAsxCv79m3NYXsD+BExL0XK3QKyzgJXpk9TXbyHUv
wbna9ITkEipW4vKXbC5UqQpW19vRDMbNBDxtCZFhdYJFqfy4w1XMCyxKjpefCcYN2M0FzvbOQlp+
qXIV6AiPgvjb5LNfsO4kvOKYKhhd5LXRupm8Uu9q3HMDbzsZHACSW+Auks5a8qo8Aoldy4GHstYq
laSkB+6TONg6TwLqiBbNPWFL9CMwJKdCP73vvxI4Wp1tLFG3qQeZblaiL/7bdg3ZXVYpH71e1qq2
+4+Msx8DDvpm59KDTe5WzJv0rxJ5ZTyESsNXz8KRdYLNF32zmyQxLy0nVX6SbmZhexbmqrZVBTMb
lnRpZQ2J8MC8b/JZSNf7qC1si2QkD2U/cUsp70zXEioymlRYXfGDv+VQMpCvexWb4/Q3dbOCXYna
s/mghY6QfKX/KJM62pE4L1UQ12Lu7JhOmBNUZ1Thl3VyKhyE/HWkK6X6h7NiImKOAWOw/XhruOEa
4AewmuCIbiT0H41WcV/4a6XOUK5asLwntmc/ceyvnvWhZpqSZZz2tlTMqw70IKi9Jp/jgOARQzFT
kvMrlTiYQPPZfZP6Rp/HfV5VDQppFNB6CZ4j0vaOfKbYHINiJso0NkzJaP617W26prHEPSS0bU7y
T7d7qQ9Yr5Omp9/pPlCdPAbtlAsLOKsLs02QDuz5uZrs4FrrBjybjuK86ujFZQ+fGLGg+3x3oSoz
6PaH+seasuLH0kKagvsY+go91S+EjhT8j+HlbX1nzAJSluJZC5FOHZOt7XH2t+80pwfQfEDI6yOR
XUigU2k8XQQ1Zs8/WOF3X64N9Q9URmPU0OtwXMkUy42qjT4buis4o5v6jcoXALNx7oP8B4t+RjMq
s1FrAskNd0rcHPBjOFFLUg/y94z/SBsewdc+hVQFlYFqGTnxpYFH7zZKaA6HTxkDDxrDj0wzke4I
HcZniyMV7HKdiNbHvh0dWjfnt+37XrlUAcaClUSNcQ14wTn7/RaCYAfuH5n/Y6UFNRE6L1y29k9i
ytV0rXz3nmYsnTWjkgLM2wTedVbGKHzdsLyfklm4fYNMYepKAOyrKZBwmxCokDw+9NSI+hORf3I/
FgDOrTj6ttyheDwyVi3dePmvAuquaMzkSNl7JXjZ5QUVxeqKwLAwFQLH5BC9R09n2UB8CUGn+eAe
eDW3ivsHq1UajBmqttQgntQKzNbygW1rRKJswx2to0zCZAkkPfSiJ9cgmYwVpN/Uahz5clAgh6mL
BFxUAewwx/B454gweM5oARXloKbz26ST5Mo73JRiDWmMY1cVdvR+TDvmpGBNRiforWkyuhxY43IE
HSZY7FHJkDoTIwxzDlgiqDRJ1Zfyv9ZG2xGcTEVfK0HZaBbEHn7bkkWL71SELk4v6acsQu0w6R22
vdEwjq9HwuPHs9BZOaFxujPCWEK0RD0qMM9djdgUzsCE2pCSFwpkaBBfeBgJ3uxxrJzw8NAmQwgt
RaeaTf6ItxDulrAaDd9J5qRKp8REccvTmb93+94pIiWJTxJd8n/r/BhjxgW9FEB6Q9WhYFRSxYRV
Jot+/YYW6hFK9h6VAgyM0AU4uzU/F5PYeSwS1JD5qfz0hKoHKyH9ykqj7tDhGaXcY23PvCPoNuCq
0geJHRheZv546kQPjjCrI5JXkQaieenecO7E+lUlVcAeYgF2PK9VpN/BYGcJJRMCIihwP+M7/mu9
1QPPD4m16djsYmQarCH2dx8InX3BGdlPeKgJPFyZ91BkYOhzEs9VAJvLBCQmsa4AudOQuV1ldFhV
DbifVHtUQXM0VJ6RkHNbKtO3zTI3CXoo9irE6sY5AhOzm9QSM8c5l+i6AVdQ3MtSJ+Ei7rWcDkh9
9eJuskoCDvKFdbbqZgPm14lxVnwoPhKQ+lziQeaCYwWDD1BBFvVleXzLeLJq1h0kYFk1qWXkchuj
r5K38GjxWevFaD+a2j2mnA7aG/XCs/hJgY8wvjvWiSM+GWHtKOZVZJs8qRE9zxVj5x4brFeALmhS
h6vtGErIgqhskd7PxyeNcDM1Qnfm6QAYNuDLxu22fdkQ/4UtoRMq3ECqL9iApCn01n14WOBF2N1I
MhX5Z2OLx3DOhidmDTtZIm411KAJK9iRb+3O1bSLPrzgdEZMMLJ/XRuoahq6+8JL+czzL/PjIHJU
Rje4Fho1OGBVHgUQS9DcPgdaSZ9KF2Tv1LzthDGq3K9YFCbNYdcCoXU+x1tqeenq22uLIy7EYcQg
Upu9sHpuasqjS0MnNi2+dvPonAlFRHNdBSwMMj0wecP5SzWwZJkdmO4Wis0tqKCY5oASg1eAdiHg
ICWumuJWkALld8+9KjUNJMNavRjg3X0FBuEZFciVR71EDRaNHR1o8LuN7m7SIIHOG3uYTZ//0b6K
oS0BmHpmh+wKJVeZn45ifXMsaAFxt0Yvzyq87AF97iZ0NvubSElNtb2G2nToFfupfSSsdGfH7LFw
/+3V7YtQujfsyRdK6gywVbWT6JC+FVmMTGNp+hmNFW2ZD7RTeCems5KWhDrLbLuyf7W2TOkEcX6X
zPQjpOB0P+f/TlxJeDmlWBGdAVBUOy37F5DkJnxYlntGJq0MY20V+BQMuBtvhsEqwfUXfc1zbEWa
72IS2jialKa/bbNlhWewl4e42Z6l/L3VIdnlp8jGoiwHqf9bha28W/uJIKQl/oZ5AToupQC0Zue9
9ERQYJSYn8g/t1mvNnW/SNNLugdY2kIweeY0kvmFnRn+ujoGrAxyXYInVp2G/jWUIXvzblt23BaV
bceM0YyNgiEJ6wouDe+0n4tyRctSImfegJp3hxcgMu0xxnv52IbAmiNxd6aibCQ7lCsmQbHEaWC7
Yew8G0rI2XnFd8fvkTTcIGfFz2idhaO8DXfs7OJ7qJZxbcH8No92bKVrZq70PzJrpko++4PgWlWS
nCZzHGb6VIduJ6j2Wjc5Z5TZ0Kr0woGTdt56ho7i109rgl6r63qvhdI7zaXM48reIElUrdEV3DQ7
C/h1+Hba6ghS3cnKcLNEIrOi3ihAwunhCDXd606+7WOuqwLhJmhFMM7RlV9qyhA74ytotVBpU/cJ
XML+q/eR7OlGHfgAOiuDhY4xQPIM9h81s6sjColDb4oNjbqQx35NejlqJMm9Dt1gVF0U/N9ZX54f
nLk1uPscOX9ENAnLjXgfvA6DdxifKRyLHjxK4sHM3pDtrZWMmxP7S7ss6kqYfOKsd3izAj3E3NMq
Fx6yqaj3AL6hr5P/VYSmA0ZI1sdy6S7/+YJtx18B0LlGjivTonl4z/m0gUcuXDlbIZqXJ3BCr6tG
5uSiEeAX+KrhltsBB5CnoJv0Zi3KuZyJb1zeI3sF29wcwfK7qV/NX8nbx8xLptW7Pafgsgy1DxS3
Z6pIIh8ISah4JQrSnxfRlIoqmv+XqeyQaU1H7HWf5NxxlZ8ZYJxV/vhvuEwNb+iWdTPsm2PqAqZl
Br+vbMOTlQU1h6fShZcdD8IE4HcLMCNYdmYQo2K8SKRjrgLGQqcxcpEVBJwoqd+hdQhKbETSuVhH
znW0JpkZyy5y0L8+4h+OzBfSTF7PckSnu28o51ROpI0vLEm5ZHf/sg8KL9Qfuxe3ySmLH7fiTxvY
qEMF1o570LU9P1i3geDQiLnT1aPwqPUo8ciZDDwsHsSz4PvYvevSIkLXK9ljvdMK1si9IUPQGaI9
NlNsKgW9zeku0sOvqqGMIxm23nw7FdD2ZuyfTllG3xKq2311hx50eLFEgkWEC1GGnZFtOGlsKUbp
+pzpvtAdczIrAFR2eBvc49BWriYxu4W5WtEWwhg8So1bD2btmanSojinO/oTAEDP2Uy6Lixo2R35
tf3lGqbQ3HX0pseh1cDBD9EYPjSbTA2o9p+GtqEPod198Gcg/jd1q+jjz3ZVh7T2no8OXvQScfNp
CnOFRQFNZAcpp4t7wt/dJaYHzKjMnFxqicnmU+kf5OKnvs1HhYp0uK4/CB9+J0E+568x9830+qbq
XhjdEDViTGZyKlbaSRV+TY+Dtk6hOy7Ds7JKKGvv2m0v96F+TP83Yx9UzIuAFb4NEYl2JJle7WcZ
/00uyvT3SDu9laNjhs2UscMVuPJHOXvIAoHbz0tmJO8CvCF0uG/PImGeLgXHW1qOE0TlK1IHtOoL
bRqESfJywhdNafmW3FTfX7A5PYOIJbaK/tWH9WaytAwkt0zX/yMzNTU/fPMDs7VnU9i6dwXxS1jf
KFxggUXGDgH1Slj0QafV3vRq5F3S3cWwB6AHN9KHkziOTUFkuGvoqJVyFMDh6rv1QmhTXilAmqHC
+ai8c5LMDAjRdWEKKQOW/4CEigrj75NHc+ikFxtxaQu42rjfxtIXToY7d3m2a6wG/DWKl/hx4ji1
kY1rnp6Cfm1LoxwOiQbbDypyp0ymh4WjtwhLh/f5jaIh4u3PcEUwC/BtZbSKnDvElEfb8OuyH7O7
xyAXRLQb0poH0dV2LimSsjZpV6dsEzTdgcBrE+1GSC+mISNN3pJ9LkT0Z3bm9qE3kSXFtbyj9Sl0
N1hdaCy3DrXm4fj77UpGC25kyDnAl/EoWCAT5tsR3Q2b+AyAd5ekChOTlwHMjPdwzkXTwoNCFZ78
C+Z8X93fqeGCkgqBMk/U+plob2RbXy90XRb63tkjtu30uGwpgxo1NT4ibkYyrX19ct2VhMBmbSo2
qvisG1Po3pV2KVvniVJ1ARcsP7a16u1AjDB2lmLeEV7w6wURlAGbIyVMCwzjlaIGDvBNVXGahjOV
lbth+OIJNjBKUZyVvdqUxFGbkZ2QQqtrTFLZxh7r04iDDBDvM5NQEHdKmYMKi97DmmwdZ3mCC8kd
PZJD+NWppEXhzmyQzacPiEQg/QuHVfI47QVf+Ayb2ZzPc+vMjQzjybXg0RY9j33iU0iI9X8djHsw
z71mj++P4Kan0Xb0oX1g4LfcVHaZ8g2V/MpSYu677S3E/j4Z2VlC6rrPpWVqkgj8/8Q2nHnOq26R
NjwO3DxOzrW6Kt1OEdt2rf2GGmgs+GVo9Lh0cpUL7xdKuUjaOEQGLR8rISfFlDB7Mbn5jnrxYHRz
ORCzic2O35DfaZd1VWyVIBBKkqlxMnFIVoRubYk6U8hfVKTcmtOpS+1OdDDqYGIgzN9rKzRD7Ny4
JXjuQ2FSCDurrjpSz57zuVg/8aGDTn18OSWu/cVcSjgY6CBJws0hVusPn9VThJUgzKWnr8fJ50Kn
ji4rMOKOziMi2hpVHtqFnlX1zCgpVEMqSBcRZ8Y8tOKvI90X74kL0a02yXip9jVAyzTZtRxjqj7n
39lmMlE5tSlRfBamcf6YMSjLvOAQFAG3kBg5MCez1fldVYQucng9+SG3l6JcQfd3W1r1zkTagR92
ZKKaogCss49UvTFE1SbmmyGGieD5O8WXQAOwxbZ/eZgRCdjXuBIxnoET56HDhF7t4gr1sU7a+xl5
vpCq+Ci3pcxBjYVVN6hHJUOA3bvXfyDxSwyfQPugrjGSL1R9iEdczwuEIooKvqmDYJp0iWhUmKaM
arY3lQntVPFjvA8r9q1G6J39Bi/YoSP+UStS0mF/i4FGTjyo1rqZ9ouEDd3r17gwx8DSZhkz9h5Y
Q5sxmeBgHfXo8ga9COH91MFFMT+yY3PbDq6fQ0/oKTBKTSSSTDWSME16fHVcDoZKLdNgZ8B6cNMc
BCeOc/5rQ6yn7Fb8iXYY8VCDcYkxSkh+QaziZgUzXb0bQesoTML0+8LhjSKH+M+7IXjwp9UGRNNS
gbJWPn/umIQEttqEuDct3FxLFq3JawpHl2ct6c3gi+D+8kKrV5sfB3N4jLWAZM0PvHa2MO0qO3hV
3UrHrrPJhQHTjI1AfRsONVP5DSKfisoJhPncukqQ8QYLVVtpM0VFY9mkkkwiJjyHqnx3F7m5fhgS
Xu3c8UWPAw50dsNLDIDzaJCKywENjeILebAACZQ0yNzGz50L7ExcsGRMp5fINFLJUVfg/KJPC5Ib
i7mCUeIGFRDh0KuFZ6vihymfEC83WIjNRRFxnhKZr9u6qpuRe/epO+oeZd5CNiBWfpke11ppFwmK
OgRgH5UjFq8Mffp7lAjBdWTDYgbc3AkdLnTctWjK9ppf0HcMtZFkYenZ1Q0piNbJVWLbduSlLeuE
T3VptdFuC6L7Lb0S0o1DPbE5h2AsoWOk3nFF9ceRoLs5mMW2eWiB+rQJAdXuanTg36t7BNj2KdTV
O4lcrDWy/XMCqqIprUYJ8Y/GztXFd/dvP/umnc/KKbax7U3jysmQkJYMGSbSlBiKQwxzHz57Ziqe
Fp9qai4Uyinn6iZEHV+wdvVtwvkePElJGDTAFukizTNsS5AssnJuwM1D63cqAMnEjA+DiH7E4Wo/
l2n5+NByUG5FEyS/4b3/6j0Br4IoEcvuW5i/uFAHEG7lqJUA/oz+dF+aLdYI2DoVB90N/4RVhkYf
DfHqzU1bti8eUECL9B+uNmrklB+Z1hQcPsxYU6lktwsQHuI4avxacwKyXwZoXaHp1BAU5Vph2huJ
VLfRKQM30Q7cm8R29S9ne/0/+nZBX/IQXu1VlFSdfEjDudF6ypAtitzMLth6xJgzIREWlPgG8Rn9
6PfHmFKNfCVBNtijunSkL9wR+P8Lo2UpFMDPtHzY9OMSS9TSbxTEUccIXNIoXz/QsyJrt4vwBTd6
nMDNIGjbi0rw54oXKC7unJGfZe6EpAEdqZ3sK53Uyh3AamyBSCMv4+AeTs8GHnyIDgjyy6aZHqG7
+eTknA641HWlRF4VJ0MGjlGs814slXP+bVgZxsac5jDhG+XgPHWggdoBEQkPKXPbqkWrBx0rzDTe
ZjYWguocikceZpnGyqhSIizPQjSCHYKXlT7KO4Oy6JGcDUI4WR0JaByaNdB7SXLrX+Jq9HMH3cR3
6WpfMSa980WFg35UIAQ511hFrd58LaofzOlY6fHqOQkia3U+9qsCk1UB3Jnbs0ny/pr0YcldHQAc
BH66ocQW/ioHluM1Iv9FPXpwDoHc2OwNMWLrKBrTVya38rTbhPtgQ0F8VDK/RPPNdyUxfjXOi9gA
GgxB541mERJCADDu5vc/jp9CL897u+3eaaNzyvkcNfldao9VI1ziSvdXuwdEbdbjI/KplpUouSXP
5DdNAbDMAlW8dLUx7LejL5PnIlR/ptfXxlHIJE5JKqSGbDfwXQDdH5uSnlP8y2zh06m275Q9ty6x
LDq+b9xuLL2kLUB0FBcz+5q3Rak/n1nSRImy3C4vwm2pndYth+QjkPYJedTDiw9zJ2EKpQd099Dy
h0e23hpANlDtRYtgmfOa+JDQIW9iy10u4dFmUf+iirnetSCPmBnOHwkXZXXEImkANFu9xGZAKUVF
gjHAfGL/nLgDLjfsg+u1iC7AUxp0Z3k/7StApMUQ+gGTaW/rA36RQGl4kugJ3ND80CiOrfdb2eM6
T892o9RmbSr4/Q7ab/JN9AeDnxVcRXP3j8mTxLdNFt8Enu9RieZMAhHZ1e5SYHmNiSoZcrDefLbY
j3oFS73A1Q+jnu4vZywgibTUf6t7NchWXegeFlNqeGo+/JCG85LGnfYGg8dYr4+GnFjmvZOZ+/S6
iILd8PjHTFbFaBLumZuSr04AfrCZ1sZIWFKr2DvZnMKS3mxZ8dtGMedJGyqPSH6fzvj74qDJO3Rn
JCdgwJvqNEknqyokODIrbLg70EdtPej3O+vXK1Urovxv31G2uHlA0ZbSWCF9oYyYcHBJVHYd1vKo
x8CC+FzyqhaDUtdKWnv+hYfiH/3Aa8eK4WoqHwleeSvKYndCCUy90ncDVF4cCywYH/XsBtjjEsbS
Y5IPmYM9sn6dbWQdr3rEPJTJjo84kojJcbEqFQMfh0lkHKaYO+MPR65Oy9fwRhOJGkyE7u8w6yXW
TK9+YGfQms0vhCcIlvCRvUsXknlODnmYCJszWi0FxXcy4ArAVh0+Ld0UNTlMuOFTA5ll0sCbq76c
UqYqxINf2ZAhFovluEW6P2TF3XDfffTyrWkoGf8n/j9aT/rJcGPvZ4ARISRNNYqizOJobd/2RrS9
XJ7fAAdXP5bzXGef3Ls909TLVvG6kLZxq1T68MlCp4lsbg7/B9SLeotXKm//GRPIqXJFg+syKks+
xNl0ZwvEVGxxtw43zXu6CfcsdVRKdWnnqfpPxnoPqj5HkyrXkixO883rF33MFyCjrw4fE3ZNOx/S
r7SOBQNBsooIXAwaupoNxeWzFjDWF8yAn1aLSh+9c05kM1Tw5IspbVfWXRq0FAt3cFsaUiKH8ELD
aNrAvQYlb+dnAOO2t3sAwCgsouoFD8fJfFmg6gjEErynTL0GPg0P9YzJacGYAgnH7mj8dpCII8lO
/dkvUgNdfzwlCoF+l1CxNwZ/5t+8o9uCF0NfkXATCHUDBg1Wj+65S8RmhVHthceW7j1gggMqKVkU
cirTGcF92RV9pHBb5tuSuY47206+urPp1Qij7olOHS0BquleroeOjbFE8wTGt2DZDBbo8DfKejNj
WpG/pKEUWdm+jj/9vUGXB9/uIjN8fABVy9ohE4JcGJPd/O2+H1cPYDGkYIdOOx2vS1D+o61lfsfH
q1XVJud7tTbdZm2iP9nRDQkqtA/2lx0vWjI/KffPbBwo7UtIYFXzk6sZ+JNud0Wz2TR6w9nzgC0X
LKtQ4dfjEKSUsTBErjwL41w/DoPo70KCOwQvCzXWvAgJxEe8QmsfAmuo2AfzaUCkiEe98LADsSHY
Th7bivt7WSz6kguCO1tyJnRHHpyJj+q5LP/nyDxFk2W8/BePPZgy/zNmXe1OG9JUl0/UQTKEbIO0
DYNF97FvW9D3F43NB9TPCx+DEARyXTQMOVsEr6MHUIMLOrFYsr7x7pWtbqNbl1m1FqXpRBOHM6bD
ejdFUmp3e+vty3I96MpBpCuH6liYlg7qAhASVykYoJpEqjPcSiwtUoiXXf/44rd16S6KLOW5juoH
aBcC8V/82euMrsehyIZOxRnexOtFNns+yrW2C7J/QSIPTSc5fi+2ZbHTPD9YaYA/GK/QK/DI3pOf
tct5jf5Wz/Zmb6Cc5T9cvG9KBu3tKaaXkPNa7Q3TDfnV3/w+iCDbnuIRsxwn6nNM5ecKyGwc+VWK
1tVn+zXIVPCwsgl8kwIlK22UfzIXimj+yJSOAQSMAgrpMNm3Xj0wX9iZCZDGP/t/jeKsZLQyaCJt
xlspXUGOtHx1zE3sFEcPC1LmT6Pndqdm0dUTxxjGfo9TTtafs/UkAM/ig770w2cPO1UsU+yJTwH4
kCbSeOzHiZE9xD80tJNAuY1Ehixo8itFk55M0q+HOkYhRuJd/L5R/9K7eoE+vjajbFIgcdE5rWS3
l9LxtmRGn+O5bW0qY9RDMMyCfBObIMiKiLbrGNQzXrc1G6QRT/nFtYdiCkvQ4pdgvDcRqJhJDJZT
tZoqfhPddY/ogplTj2ZKEc8A9J3Jgx8r7eFwEPHW7YCl6AVPg1sGpZlkVOmkn9vSX93IUJ5qI1+5
NW/CmJ+kLufQEAQYh787UT/z5zTPI41Uj3IKKo/jvRLUGRadYDt4/wudZPWACW51Z93lpYmVh7+s
YcoZ5tOig0/bIr8bZo1uKxCakS1jKXLeiKPE2hmXS1jD3HdKerFpvg7xNjHCeeU5N2c8id8r916V
BjQESlUD6utt3rbS6jYdu34Iz4FxvDWvMpASTD9amI0AqGUsUeDUmAce6K7HeojD0+/LJHeIWJk4
ubL+AMc+CfxA2HMKPeHp6llfrQtj6BC0laW2VgipyrCJyNq6nApkdGha1YE/9loG9xM9zwHq/Q/n
6WeDEGbX/ZAjdyA274NIbmDl/Vr/xjp87L6ChS9AKM0W4UEchbxq2xjPsk4iB05FU//r7MKIIdUl
5RJRDPw3P+GlAliMsAJYxRL+k9JWKLqu0/Ixqa88HGJDv8yqVgC5qqPK2NE+mSVVrw0/ecCGZx3e
B0z2ih9X3SUb59PCqfQKkjzg5yP2Nbu4zuPcqhSqNYHJHkRaHAt2+nFrzZhwtW7qnmFOPz661b+d
COuuD86bTiCg3uxJfZ5BaE7Uo0eL90q0jzAl5io2gx2I568okjnIn6Z+AefGRVNmlI1VWCM0u4u4
b8iy49Fci1xggSiZfkZ+IoPdQTbEZMiERSOPUiPbTCVtihbrDs9ot1kJdLYXSS7hmgLAcUDbh5Ce
sa2xk3YoGS+rKONYTfaeD9JQQw9N6w7D8cqIdeBWNuXHzP/bSxuT+fAzCf5M9RHdM0bsho53WCFB
3Nxn6eBqBqEAc6x/C5DGpG279hGspdLCRJ7xN55EB/DXoKzNzoV/u6OzLIuwSo37Mp4EYf47zzxI
4DOn2BNLWmY/ykiNAnnJS9S6bVHEQqNgiqd1MUl3d1rHzu2S7VpOvKOAWW9QluzRXkX041PPRHfg
g9jhXAua1i/go0tKMRDG+Zkh+IxjOADAu7iNVcj/nM5s4OPEdaWMFUekuO9/9cEO1lWNb8q3uukE
aiibAbYYOIX9LGTlaZjMjAX9VHUcylClFtwK8V45Irs+y4ds9fvyl3RYf1TFHog2ii8Nfuom40LC
eey5y7fVC/505RjLfxVcx2TcVOk/Im6/lH9e8zLsOLRomYfsrhK8NwWuE1fwvfhmH+YW/HuqESxV
BPJRQMQbn3ykgh7w7JQ4inT0fFlHaKDkpHG8TDCYF4tRt5mODS9RmT2tlKNBwjwwPLw5r+fdefJ9
0HI70bCNW8Us3nSAO3VPLQbI7cnhAVtM2iWAe7kBezBQTK1sgYEH5sUiLblerR3e92LA9ADNpArT
8P7/LpxlPcrgBgaRQyw9KblEg0Vack6rq9AJKmlHowCrIpAbEx41S1a31TPEjH+ChnSWK5zvT6ED
qfsL6fHDznTOYN7CVeh8leTbl2nu+nzDulK/qucllviOhtw8eMdHbF1H4XpysSTO0kJoALo8BudG
fj4zVKRPm+o8wSCZNY+iELrKV88MgJ7EMPjlguiynXmwwd2zcm/VcbUjFwUkT6+A3ZYAqIpS0rFa
8bydyohAq4bJoSAaMiHUIntMeorLHuQd7zMehwPlMbrhL7slZ021OjM5m4gt0Z6pKwgCwZ7zITnT
ULL14XStKSaiCfAl2xR5/7i39RdFox1/rbAMbzmGXnBPAH0CQ9qUkSeGsFsxWoFwxdSg19c8gvR1
CiCW6Eqr5JZuJlJfue1hevmC6nwTR/wYXmKm/STYpOP3uJKMoGXvZBHka/QmvGQRFKXkVIernFf7
AnX4m5cVNNF45tF6kdqfT1O+1kisPtEkqlZX2FiKAIPABwjhQwehVEe9mMV0LEwO8XZp2tq1PMi5
MOe1W4b45jL9O2UO+F6QlCM7OWCjabVMj7DSEwGZyKNO0k1dRhIFSi2si+7ckYTlg1hveQGRxh1h
55LXlCULxfiPyWLP1Hc+qO6p6AtkBM2fJAHIF1bspdgBChdGBThhA/qb1MxReZAN1kpcGrb5mG7F
LKscdwYNI61X/ukSjxAnXqLsu8V8D30hE+0ntmYxMNspqU2czRB9+dDnziHW0/ZeAeMM3rR/NRWl
qwz0vNP4hKhfWbMOowvzr0WBss046ONY4OJdiDnUW+ZK1YmNynxdcrNbeYVxtc7hH889762Dv6dP
WkOZaIWVtZdxVYGPLL3Tx0u3DG7TF0dS1CohoYvZtoDZRZHGO0lzhyWAnJFUESsjycH2Aa6oT4zp
g34FSGQ/EGDj7Y/W2b4puoIbCSQPB+vbKVGQ9OgnzA0Q/5m0yBezDPkv0m+Mp1G2zHDo7OkNIfza
NoemwQL240tNhQdslWUgjrePDrB5NyiyemMOHLoV6Ono5shCR9g1W6e845wYd4oHoFVh4bIkHC/1
FigCOtriEAGdZtaJmarD4t53sl6i6AoYXPsEiRbLwE6EEUVrdFQ54y0kmdIKXPJwuyWEU0edhkRG
fxzjolQip+arQMcYworasbTQK2/mZE/T33lmAJkGbrKVcbMDVfOINLC7rVTfLEPyP2BQOMiScWhW
9ivNqlJywkMyiSdrG1E1QtbHM3KHFaoPu9oH7eqokr+ELcfQi6reSzCh5YgeDzxGIFrIR5YxWRxe
VZtlkpNeoy/0x3Cqsud3JkVMBzdmwo0KD9RK3luq6Kk9tihs8ikkrk1yGKqiQWEyJKVYMuxd4TSK
BzRfmS+uhPbqNeSXHyOzdD0qLnayqoBmFz1+eAsIpB57lbk58JXntp65puUjXSExs5DYRP/8qrWL
RH0UH/S+tQyAneCGbapq+bipTM6eWv8iOA3ja+hBGmztOY+fU/RyTMsz3xMKfSNte15vbqjl6gO6
FrvGRYcdBP6dlZiGjHah43QmckfccrIf0qBUzNg2Txyw0224zpaASRCsjAgAjwcICB5YavKyeVMh
KjvMEB+/HTSgbQgtrJeYBA5w5ZpEBugyDBJCHxQz/r0p/5laDS9cSca5pQvZrvus9dFDua3MYZp7
tGE7C9/c2flbLTIc0wcbD3QuzrZN8cudwp3enG+g2ceGgv09NbjFhw69+dGT1E/SBYUH9NpqVFlw
hjcjw6PgcTs+zMXuTaS7brfPRDtDt272NZ/KxMnKqKMiChrJa83tmgs9zXlnJOHp1GNzJ/KAWw/C
3ZJC3bYlZJYs6D5fJQ35G+mW0sCSCAnjSgZVc6/6qQVj4rfcj1PzwUP2hVjK1MY6qxSwgzm/VY91
M1Jjc/3V4ypsIubBAXPVVgcgE7MeFd6EK6A+5CtM9ewx70gpzO6IAPZB/SFj1/6t81G6iMSFKrCk
Pg+otEtrrgnUeeM1j5bHC0roZv3JWaRL23tIGBdmuIvFOO1b9YMvMLgH/KQyqFiM4sIcQvhKVtdM
hmKLCHdK9fwLyJPtwCm0rRukfJ3fQlMMjRZUY0uotUrTWASZTG8ctgpAE2C7C9RBSM/KjX17uezJ
y5pIQ1F0debg4CGRd8CoCXcUeIpFgGGVtdv1nmfkQxb4dMbym32dZ3jI76rzbENu833HmTQ11RR9
EhmBzKhZKYQtrL/fMZaiYVGlBze+xGq89TQZO2nZ91EcqvM81NVuKpirZrpJezKIEiDxwgk2dUrg
1JE+4dJ9BbKOrtjYfwALd95UhQ4c16fqG2MhlBOeq3aFJiHYTYYsaTB6eNAYAmKpGCe3Hj8iwjoN
oRfK/mF2Ry5ef1zMhvM/UVCh/dua5TwUb2ru2n9u2sN/ucJ0nYa4SIKhrSpVL3QaslMoAvwK7nxy
ljjyHqvWmX8NG6/hpDZMQ7xyTF1sKoBhF78yejnIw2MCR3d0rAhEfVqJ+NOMK55EcEsD8SKq/c7F
6+yq87b54+pF2IOloiE6LN8wSzRQSUpA33jyoSm0eJTDlviWzvs2BdTjT85gjhDTeawje5IZxS66
8zaP00KDtq5/UMtHKDL1mDuk+8+F9sPCq28mlZFnJeX5GkRVrCVTebaGAFZT8tRD04LzOr90xnBl
PeuAT/6ilG0lt15LLfLGHS0ZMKj4+ml1Sr5ZNj4YYqkrrYXk6S2wbLMgOPYBfP5D4dgemWxWvSor
t7C+Tm9zelpKnqsIw7J6TGxgYVacBmhgXiM/T7LY3tnE/Y6FLnP7CK2Leriol9BGuklWlD4Pv4x5
/4TnGxVy8VmQCdoG8CZUpd88ZquGXjjO8uDchAqh/nzg5paF4QP4FvzR+8Kdg4gv7SunAUuwv6t9
1uGr/ZnIZIG8l58OazGfllCY2IpphszpmWatujNjALd3O3679yYvVbuGH7kdEMZ10L8ziNWFDQkC
b1F5qBF6FiTMg9w9a+HJo/DAYHd0IHDOGajgX1d/fe3mMjXMrWKDjMGjLWQ3CFQQBlQIre5menQt
IozSRr+dhZO89oeibeF6AGoNgjYT3GuRYtbH9+6sgnxnL8s4y5wH2AbqOaovv8uEbrpA4xThzqyX
qIYbQ0buZ/l9ALfq6/snwcOVxbObwyfh2bQgGxgp9ToFAEw2LiWxCGs0aImNcaayWuL1oMvpccOe
zd/XD83V215wkdMiCD3ol/0+PxKZ8sjYjqm8DgINB0dPbRpXRIPzHLX5yFto99iJ5bGD7GNIaLEY
hrK4+8mb2NhxAY7lbaA8v7nYKVL3wtQkT3SKW/0RqOp0XTABgr6gyP552xKxiMsQTHBHMT4C8skv
XRXSFbibkmPrZyw30IzNTG0wA43WHLvCTKQzIcaSLV4VHUcY/Hwq3nze04ZeR2vMkCNLr7yNPoLx
8B20z9J15bXOTKzEbLiGD/2HjfipFWyltSqZJPFgGcOWlT5JCyeKI5PHPfjvCb+t7FTt/jrKPq93
eUyPIO7hrkNJCOdr8P+M9gczyy0xbVfKcFAGwp6JhvsFJrjF6aEdsC1gBo+AiDG3Ow1C9L9bNghZ
um4NEfHVmlfsLRbKnpM7CiJ2F/MZa39Pb8eRc+b8D7kumlAND6YVzHCCkRUI5ga3DC1chFpEYaEl
KGpyzLvJ/9Hx1ogS5K0Dr/bE+cwh2+a+H4FGRRNcW4H6jX96u1YcSZUmLcY1RiN7qK+jMJV6DfG1
vs7vELQVBBbaFhXdAk11EKIrTy8tyHxbxAfl6k2jXC3KVcTL5UNGInSW/8OTtjfHO384+9Do/ug6
GUZ7eSp4KVKAh3+c5OsOHRXUN2uDQXT7z+ps4Rp/HokCP0BLmg0AtPcW71Vz+a8Cl7FTVCI+s6if
4BL5vZDqsxAvRA39HWiKWkmjhNErFuL8/6hZSHYIcGdKDslswJsHJDXzSvMp9Xq5yzhHpcY+WRqH
QcF0+sI9+fGI35Idz+p3feCrNGclzWj/3r1pbQ7xCpwvnIOFjueB9N0hgAm8Y2XD9rEFBbbBY3j8
2JKuZWddxq2xvwEz2iZvCrf99pAmRuBsI7uHwfKJKAflmjCeYlIo7lMUk8d60Owk5hTnQVPWB/LI
hrME3/IWLNxD+QFG05KgtCUC+o5TbVneCFiww6VfBMhiqFp7lj42a8iIsv875HzS4HtOKV7eQeB3
kYR4jXm+kqaDjUTM8IfE09rdMu6V8Wq9q6SqMlhAz7pSO+6UY8KlojGuG6upMXNbc/V+ouidBSZB
x9wiC/1fLM+h/ChPXBnPkXkGh9/ed3FbUhCPm8oLYO6NqaJ50haUAdSBeUOppZM+i0rOQME3e93b
g0Jil2mS+Lhqn1YZJf3KT5zDyitjOSqvVno8UfHWYaqd405t1IFVgCuldxLeQXgiXojd00VWyTaT
mFFKRe4l/rs4zebfKt4eEac6rTmdd9xJd+OR1P9lI9ozFmV5YIRXxxLJwt7ZmplYQbS+S6nmpKN7
3/iqinxbGWt3pBuV2CtK0DU31EYcUF3Dg5SFh7nkHOu1wjuqPKxz3x0GA8oKUsfhq0Wq9WHDRfIW
615MLWNE+V04h3gqtoF2Qxc4vzTENyRSREuDBRZYoX1WlHoKDlIaJnQEVWVnnnbEagCIQJvL9P0k
hy0/HzJB5BZl7uOeZcDahs4O5ncsTZrxFqOLx9TcAziPdaw2b9Ugp4GH/Uked1RcOyHnXPvD4Cno
KwZZ5zCpqNSlZnv2YTGqcZNkJRaZcgt9FWzDydS7H3rU9C29DPR1xQP6BVhCzth6O5vDcFX34sPU
IEprb7+G2iOJXRK6lltlBbuBa/+3IXagkfZXIkHjOlDdP1xS8pGSQZNyHG8kdH9wUc/UJirrfamS
dCIkw0k6iFqwfF/D6KF9K+kGL7jICRuWTLBFjGly9yhWcbJ8vTN5vXXACmx16WLa9x6j9j2/AZyi
8Lt8uX0teuuluxjJUsRcp6Jk7lzvKtPZ4ZvLo+RHnIsxjp0cIlNRgE7xR9QZPy1HyAdDTkMKQpWS
PWgqX3MUvpZKlvgMnSM+op1gDh8h5Vp1gNgEzSx/o6wyCnnSUWEyMnKk+BjGOrHtXvqE5pL53mx3
5uO8gLd55P2DPC0ocLIuzo4+Ts5h8+nGX8C2XRigwe9Fb1RqcVlI6zqzeuDnqGWtRgxOSWdWu+vb
MQQc37j94pJmrwUvZjE0ydRyszHemsFpZPj/B+5pR9vVLqTWE/EG+AeMhlvy9Y4vi0snCzsHDvzN
FBK68a+MR/mFRgwqPOVmvX/PvMuDCVSEnhqKkPBScMIXTQ7pNzNMZSL7oC4Ez8btTspZBDWI9qRv
SZ9mDqB5joJYQ8jJskfMrl4TQtGWvhYzFaqBChCJxVDODmdU+xrrmH+L9vpqLb+FoN2vQSU2FYZw
Lr5dOjm1aLDjBfh/wBK+4g6aDDnDesm0XEzNwdOJrlREevlmKhEULnljkFbUk3hOOc3+ytpQerIB
UZdvb0hpqujhmwdFi1flThxwPFmDuo2/c4MmJfVmWxrEt0DITZbAg/emCCBg6dVGqNHpEub+DL8E
scP7CMjRuovHt5oUtKFZlhz1szAK/KUOsBVaKN6fSGQeFDYWdlI+6frJDMbd9IQ1B3XVAHjEfwVH
poIDWJbayKs/xIcesHmMdbaQjsBPz3uMOBqOecms7KjIAS2aM+VutPvrDHs7ZEssooI4PFdZw3y0
hQB683yi1On1OmMna+RI9zc7pdGQIw04yYcym1tEKyfDB/SA1kdEHSY+Zk2M1Byk/ZjPffJAZXPo
6meaBUGR6yIdKqY48Zog3w4sDOoRROIe4GwU7U24baufm4nfJYITnK11n6gQbHrVNgJ5LUb2M5h1
tW9twz6XRzVOLp0CrXXdu6eKGx5p32Oa4UuXSKA53I8RBbtEhkiMZ6wFVn/jMbB8RVyfR5lMBLjR
tZgJIkRljf5r9atRgmf9CnrFy4Yy/4fP/V3en1A4q9lpCETxAspDoQu8uBbznv6iFftKx7psWj9B
XJZKcuNVTzSRD/hC/+3JWT9gyEEMEjhsdS1nZqt1Hf9y0sO/ZInlqqCeWhZHpo0wVzw1GcgH50kx
5IkSPQmsvHdYCpaPNSS0z+GROyGoieFax2nWt4YuKw8Y0KizYCzYy9WA7YFDZAG0UyNVTBnOgrhZ
CS7uUPo4okXRvowcvxQAxVcvIeymqHr7OXXG2wjWZ2GxraSwCzVm74XsFNndd0b/f1ivTFGCNOqu
qucJc4chiHXrKc0m+HFnrM/gdryrLJ1m4NnlCi//oYatilKAWQon9fkcBou4l2SjmnVlBrojKAVB
nilOGZxcX7MQU3T1/jQVYWrC9t88Ne2KmRR9gE1aj2ur5HulA8D/lg9CfZazUIdD95613uWtyQ57
2mFPr6tHtMqDEegjNamIsdBqWsfnyk0mren3aAv9FRQEcWmotaCWGa5liStSi3x8gw2YewZ1GbqY
U+y46Mns+CoFAbxSUrQFZUfbHBqaL6umd9otJiqHlhmjkdVAXqIbFFUvvci0rw0rFf50eiv0D5nB
Wh1P9Qz448a2g7vl64g8mh67DNyHy21m/HfJOarwB8flZ5nbN9L7BJXXHQd1cM6+KCCiX/W/4HSs
H47zsTTHfqjfD8z8ng2uH1OTFmQsIW1fBaIc5e3dlHXr7s/hF6TMGnr6wuWv6JpbGXuSPpL/1nPl
UMyh1+cmSD+koPsb3WZ2eBiLw9C/yVAePhLNpIC4Y13leOfMsxHq5f+OzEhTuc0NlwT39mRXM0SU
/9XkupYaGzk5TA7xPV+eBlAje1nPvegZm+kFeIilpMvjTEbSHSd5OzyShfkb2vKAe4kQJfpUgRjk
rWRHJdE3dINBItLvDmBOsUP9VlmlMrIdErfUroVUgGMkxT/OAgfiPx62LrwZuTzxVQiFpvmg6B8+
Gr8HRi/zNs2w8SZNwrfL64NN8RnI4Zqn+rhju24cf0DsvycjYk7fW/oYOK80Vq0KlkfHLPiXbjvn
0/K0O8MgkGs4IpI6piK8ddSkaUMo4ZmfL2KUI+vV2M8Hld0Pbvr5X5ZVILOgNJ6+aOgGdgeG5sW9
/dF8BB8UwbTpGOx6BrPpZ25D+VNehjnX9SGmQ89qv8xZ1tPbhGDik7TR/rS7zvJJOGwliWDdQFjt
pKCvmsUVU8SZe3BEhKPSrrahT3RPYZMMnwxtzj4qbe0PD3Eka1pauPbIEfdo4K4RaDf9XnJxtCAo
4vDPykfvExUywVTSX4HOTGzuGC51J603VTk9fhQu8J8Q7rOOUO2IT7tMZzS+34K4gNlH2jVgle60
pEjzLpPtenHACRbNhivbsSCJPterEYbsiNb8tb1thkoIZJGUKMVxwHfpAAF0caCj8qjRmzbsqTpt
VdwVS4kcD5zOExKBJPmsBXqyMH2pO5TP3O95uow4SVXcO77NNFBDxpM6fehecs3X0l4OAvOuVUtE
cTRimEZkVPwfiSMvqsUnkwGEDBStbuef1MOvQBsB9Y+CrTPIRmMy//z0jbjzNeXfW9GpoHrdYlvz
6Nj5Q9MzZYcuXEG4tK852qfXtXy/PbP1otRhJOf+Au0wgueBCUtbRAfliKGIwIO0KyNvXfQT83GH
XLsPqSmn7UYMfeszvBs6xTi4N15FsabHCl5u/zK/ikWk44EuRJrtWm2KkAMcY2Nzh8ANNGDdhhRI
QmDV2Ubbbw0ZjJkWD5s7+FOWC8UqPDbCjJLNaIifTClks7udi5cOZbThy0EZ0gcmuNMQy8zKxulk
AZ2QCRDW3IRQCFvaWmdTRuP3ICTZQo5/eTrWErT42NeD/UFQm5+R18w0Mln+W1JCVntQ4/Qs09H1
swpxgwT4DEtAVUvbxSROznB7fdU5htZLPzPx68fLtUhl92K02Gk8fjQoUK+fIfPrp9TMB3mR/fJy
49oTgZn1hceAhFYK2nRRGlQEpzjQF/VQzQ1dZ66bV9vl+PY06i+/Mm3jWOvjysNpBLNg7bpCRVO+
3wUjXa/0d1znUvsg6EtjevMeXjdIlkHEBICcraE7wPiHKPWkzK32NNijFxrPos9m4Xad3rCbYG3Q
tX+qfDBizvlSnJ1NlnwKi8aYOIvZvmkoT5fSrs8t+cexbrQpnmJCnY4hq9k93yz46887v2Lm402c
ffe1sedtWot7sfEzcxlfwLO5yU/UDkFMxUXRulLoThnqblj2HPurQFzkGvA0Tof9wZBMb3NyhF2x
v86YAHgt6vnbDeuwvka69sT3fyXJNBBOPmN7TB6VsVjfBwS1twoZ928MumVISTdPMw6rraRunXXW
rmUqgcuOFpLchCRERUGc2rIjCg7upfLF7HPxXKyVmnfLxPAqF+9KG/g1NyiZ0Sg6eftU9g8qFiJC
Zqi1+XZzOZ9QvgQTZTu8Q485GF5syo7HYEP1ex4+oSioGf2FyKroSaR/sZmP4KYRt1FBDj/L+dJb
BtnuVsv79DqCokS5DkRuE4M2ZgGaSt1wSoDRRKu0t6Ln6AUP9louBscgbUyPxUVLQuyy23JOUm+q
yXst3ouRY36oHbne3dM03azgW1mFE6rcux/+u43svMeuhhwufPkXMwdxwBPoz0jO/q5x0F4KycdV
aAGOmA6LoaXT4Wz6VVts4Z2ZKi8+4mZQoMUI01KCkwAvqq709+DPw/aNIkEzicaU97tfEO+ZH2yl
p6IzBNyQJU084J4uVDxOtGzgH/MyW7qxdO5vWSlWsM1kmvY/FXbH45Ny5CqiKjq3tv2s7obi0fEJ
5F+5hLgvIlIhnjZo+f96jlW2/0cYaLht6zk2UIXy/NzIKbDkpt9ovk9dnPuTq+OHUJhFtK97YGZy
OiNK5uK38yyxssecJE8i9o/EGCy2qXPsq0TbcXdERAoAOI9DGzOoq2gyBrVVyr7Wtgz4KV4JNedG
pV2j5OGwya7LvvMoLSvkkwVtsUNyoEQGja9+RzjggDoktZ+oFixEeO7QZxKcHrEjD00d0paet5dt
SB8992zZ/vhUcZ2aDQbs7175pb6VGppPp603iEsCnnaOFjGCIto1iuWspRT5XS88qlBnDDkZy6Xg
of+xll4EYab4X0Ge8B/dHWHq5/HzsxhI/zmF+bbSUZN5xJRKRjuQxk5y1NenJlGS0O/hfwjG4wcN
eTccV7b+xqx+zWBnH35j7/I5Ja03jA+cfEIEWe8aMwRtTBPh2tsuErsF4xyTMplzHJyz1l1SpP+y
wV7kkaFwDFYuPxTKdhRZC4eloKfj/4eMRDHE7GXCEswzE07xl+KQyD2MmXQ1mdGkxjnU2bOhnvhj
bAP35gZq4Z5lsEXkzxv8GJ8U7UVmbQeA9hUMnL5bQzofbjjJxljlym2R4H39cX68NTtjRZJLn0oD
BobKp43JH2s0bqED4i9snuLVr93ZmYy1ymRCTqU3umdqcMLYFKxsGZB/m/YhkTfI0hG8+Jj2dXo9
baiZ904ymo0PH39ZkJZ8p66gJ7Idp8TLJOK371M8Vpkl5aFn13JspQgQB8Eof3tBLMXSira2I+dg
xnrPS2a+S0bAJJIJrMyJFr97A8KQ2y22jXXjgA6FdpQSHQy2EtQP6mOzYdfikZxSJ0UgK12vrAcs
MaQXngOyojIPxlN4Vq+j12T/jobt0l68HvwhBiNZ/+DlY3izuJJggQGuAJ92JYJYXSDjchTe+Z1E
2Y9sBAIUPjNrB4bj7SKuv04URyijq7Skvm5R/sgnl8zXE/SH9GUZBJs8H/QooWyECjLtfIvKemks
oyNamPqKTmYU+LF9q/Ifnpr9q60PZUHFG3cWMN9AE4R+wTxzSekD8LbZzxtSA7OQTpOnY4DuMU97
pbHB8Pu1ZFQmqWIp/NQkW6puuwtx1oGAwKNO3UmufGK/s++uThBaL9pCyl1CxHGGAIJousvrAz5G
HG6G6E33Ty9g3BOJO6rlkPK6Yd9u5fdvOI1b+g4+cC6jsf6+PScXVD8RQmv9zmB8jZK0SUj0FIir
qrl2PfynDLLGJWWhOwKQPAaXQCgWbsOKJDMujVMLMiIWMS2As5KarPUEEjCP+JziCmGnkrrSPpJc
tuXDpuyQljCMVALHdhRYcf8JqJvEUwHsmTT7DyaCj73kCIloBdMVx9jnDFAVeHAbgGIET+fCYi0/
Lq3ZReVNsZHhtZtpAwbdBZgh30OoLpneZdgzH8CBifeZ/izZpGbO2q0vwveUmqh4tyxOVmyAZx5f
u6j2qeEz4I0gb2UqkZ7C0crBNvsBwXac5HmHvpLyDQw7MT8tMev4SnQ8d8fpqIIJFFI8+bXsQ9KM
vp1eSmcsrQ/2rN9S/+6FFveu8gHHbn9Vo38hr9Pd+cuS7tNMPBwSxgpT+iu9DqDPNPBdt9YXZmJj
IyLN0lm/I1HDuugXDnc5Oz42IFVLiZoMlFXGdJD1nfztn77T7pQlWduicUwiFxFdFVAxxvl9OJyL
0gBa2bYuX1c4GlXYPJqdkq+bO16vdsLQhWsX6AEN5eVZkJP/V2GIkllBVnz2wIn+h/wAAfCBUT5j
KrqH4JTjoVsn/KC+vMDxG0wuwqXWao+TXXkBFoI7bpnJzlfovcC/Ob0tm8zjsi2EO+jQn+l9AbiS
fjtYIjKZ3mKs4DvLOeuL9b2xfHjzQs6Q3yUNRPte6jDrYqjCPFWlGDsqlWDXI38UXdmeMk3kapzf
vA3ASz02D7O4XKpaVcSt+ZOD05q3Luftj0VTHVBtKQSUWmxEXvfibbPsJXB+1IDxhySI5AYVcRjB
5cv2Q1Eq3jyERrsyvJND5sIihtW8tK/maCwa5o61cP8Ez6Cqv9MdYxYOvtiPe5WU7oGCjy4igxxQ
g0+9TsVikOcDNaPPBBN+iePZxz/08nEoggVVEemztsmlxOGuKvDSAwpvdVLFSAaS9Te2kR/P9jeA
5Z0C0IANrE5WHdqJjOkrhHGnCIbHds6l582rj7obf4KkdIqMc6sDXc7gE/ZvE+1rAg001956CmV3
258vfQfXw3OnusZWB+rC2ed7HoPXvC87CDNyyMYIC4P4YgxXBn4hl8GtDZoiYfc20V5OjGO+6Qd1
uiSwesdozogTepMuXlFCESwFUBh5HdVaAFWokZf3R44OuGBMu5t56jHYDy7Xf0nEKmGetfjjxa60
9bKTOw/whLlccxePp2Df8nYI5AeRbB6ijrZBuM2qtrl90USG7WBwwN0ZIMAAuKwQ46a+7pfZfzBy
/PYqCagXBXDoz3ZBMrJZJuOKOZilvRnlCcbMsCjKgCfd+cSJXDKlMUoDdfBGSnGdtfOfMmkhpOlz
ZjrWYgCFjgjISvbVBAGT1kV0iu/v1cTlIBUNsAvrkIqT1aYVaQ8y5o2gYE1ZKYWnBwtL4HBsNt/c
3R07OubSGpqZtRPv2aZfN9gW+bXRI4kAnpsXVS9iCTtVWUjSX9yvKPgQoyh/jJw6/ek2gJE4c/z3
etDBH2al+kcWUNzOR4np5upkmfsac1Fd5IJ9DHIcA/QxbliAZDa7k0y7E1xSX8nvCZBNEXEiuOJr
LbJVlpAZA73OuwwKFswsltGO/h5gnYKaPQLeTW1q4YZAP2prlWtrdYCuO/lu5iI8zFeOE2yFqasd
5LCgsbrHdiBaI59I4CfnM5wsc6fXkRhIu7bcoALQZygZSqOsKKVoXoUSdTqegRpTsB0M675z80mk
EyVij5N2SikZTg1TZVhSLfkL9yZ/YjlXznsCb6DOU2ZbV4nJZhgTBi7KZIwaL7B+a3hgnS7PBItn
holoJnKsPVJDiOukS9rZad1yWycq95f47UiIhzEhxFYB8VkouafJK4IdTJXdzNMJmGUb+aY0vaeA
xkwPujjtDP8DDtb8QMS/XozeU9znhGaH/s5++R89UZYO4zBS9yjalCeKq0XEcysom46geKHZTloB
N6OOpmNAJP5MXvwYo4GFRBCbxNctCXfQsVFcWAD+FkeT+h92Ym5nOPuTM1bvWh2bqnvWdetq45Zt
0nm/n115Evkwu+TwwfD+zqz+aEUEuw5vdGZshQuD8CnksO0O44HxPbgI1SOh5CUY1r/Zgx9C6XIo
B/L9ud8pygPQpMnDjtxifTsAeZmtC+X/cVr7d5Tgdtn22LWhkemIfqUDigSUzApsJ0gdyx4nhE69
Rhb+6SRZzIYeEvTmxg587Cdx8VyrVl4msum+uzvK2xzh5mFRCZkdkLWUQjRyydsS9sGOQQqacTJT
VPgYw8B7xYd1rfOPhnM1N5zfiQvJtJr6YDcfPrY3Po5l4If7EvfW1HntQSTXb9FuFPNzkFdzM8m9
BL4p2J1PPV6jAQ3K8zyla7CwqDjKHVwrALQATdpQpI5mgazb6ibr9nmgTtW10cyJEngmL17seyH+
HU5LlIeTjFABWilB9GcTqNNDOHsVk6PxFiHfViiQCbJ4Osf3MqRJ4VyOHStM0pfaJdRqAYMAbgHu
C5/d52XbJVAY52+6Lp1jt9FcProS+E+aSoTGwshYgk9hnotyQVvUKtpzLrbuhe2upjxehwyKEv3D
UceLDavYAuti5WoJ4Par6fmCLwNLvr49fGTZqL8f+8NyOMX+MD9cH51HtTkjoqsoD/AI1oPIzMWr
+mBabwx2u5RYvjjcwX0J4uDFTHJpPxjSO0iE6Jy1y+ELuANMBU0iEy1uAd7WJFliPljaovE4jl8v
kHdhlzxLrLhtIkoK/IYCPmoTWbgFxkx1Gyg0NXTC9RtyTE2DQD5CQbDBvBFUOjZ3kmEU3oRt/sYG
rezYIYD9pDBKbNEFbJgnghS4Fl5f6DV3H+6D6HQ+dpbVPTiavNUFdc6Nsh/N/YWecIb2dcHBikjP
U3S9OaXh6MsVZaxClyzD6/jQccOHBjhI7oLDMurUWSbXEnpKvraeJCcWgoU/vI/IyerXgChxT0rs
aOy6KiLhE36owS2h7mBlaUIqE7YlNVpiQDwet6A0qRTh8c1Wi7TO1qNQdpaYpkbT5sseLkln0kZh
R+mdwdivqbO0qUifa8RcnlU7opYMR9LXrlk0fLvSYZ31ihFH0pnwTgu65iHbCOpGYlmJkoVy8LeH
lpfg/LuRZY9wRx84tCb88/MbM/7TNya5V4eiJ9v3BX4g+ZdXWlgYBx3obewFkFK0TEAfIkaJHFpk
83VqCYlBxRz3viEzMYXV4ZJsbD/aKQr7LBVsR2emErlX2lBGpRVNk+O5ZhrWbK5r2WlgVd+tAjW+
59k+TeNvdw0rvxBWxglQ66JmbLAXm9aFDAMledmOgG1ifyPR0sZttzglTEGnYw6oY7CxrW7dvh+T
iNCD7T9q+4jm1iuJqdX8m2bjpAWeriaiGXjuycQlYuViiUh9r5QFm+vejngKD77y68qD8Js1f+uT
fK1neXsJGUFkniK5Mau62LoQsRp4valJxpbp7I7HF0lrAgQzIqiqbShcPynO+TuHepJzMJfUB1MG
rbxaKo+8lC8iSmu9/2TfLTgIgY2pvCmIE4NsGopHYDZeEHGXsrrV4NdwdOjeNK7u8c2mpBIEK/D3
t0wlYAT7wPwjGYG/CqUSImttPdD47P37fQWprl9/YxwtEanjmAmE42thXUKvGKgdqFe6qF6DWuj2
/L1dvQ0E2sNH+e3gUhakdLXhcOo+g0tn/yEkusHmr98xv17p0iEdmt6/yBjPUjdDxIyFycxg0nhz
c5i7db8uQY2XHxFGELCez65gNsfDxMSLEuoQ2Hvywq3U1XwfiZqqrrZ/KL9RcTYuqJuhpmQuVjjT
vIwq0OS/EMQS+ndco8tfJ+3uSQRqC7AiR4EPvaXSGbwPKXa5Tu0GIRO5jgHUJgrKSqWvygEeThgC
0Feg3ywP7WN+E/pxBbzNCZDDsbKmSzEhqz2I+3RhUHuEWvd297qUGZtftOy6XRz4KMJILLW8yyb9
0jcBYAgNcPSPcberzb6xKauWJ4gOxLDLCGGNGqtsD+JiHhcWIYwWlSOxfX5zt6GwZ0Mz8o1fXxoW
7ucKzORUERlT9R8G8Rp8Scc2qLuY4wHoQYRFEFx5+6nVdt4kYn2qg82r7Up3Pu5iZ63rKFg6xNq6
eOLl+2saqRthhJb940/8bhy7SUO9Qxgfj72a5AC0MVa2eaTFTkg3p7ZXXk2B13oFKp+ottcmc5yG
TpWtXckh48iY72eTqj88FMgZVYI2DdZITWEp8fPdCrDbQRcLIK5CUvtvoSi5rfwXHT96dQ5fRtGv
OW/OBLhu6BREMxZsK10Q/4/gdx3sVpuvsHyjKxOj2KEpe505h8jeKZzOG5+7Aa2Ik9qS3yFSPMBv
Flv7UGlT3AaxsHGgsZGyNXmb7ccusI3rNEoEKM8N37y+6p6haigGH9kwAWJEKNtg33b0yDkk0FiA
DK+dphxz2k/Y6HcM8hRpqLn9tDmfrmzzeENLgKVzJY6kT7ZAplNQuDQBX9IAn3bY1S0cG6VgIrAz
gD8QMpnoCwRBEv51PSI5Amim1jR60M1lSqOBtmNV0GxSzf0/jWxjCBn4LzaOmMYGOouRKfxXk5An
L8QpuHLM9/0cVJ7IkhgoxAmyyqS3h8Kfuld/a8du+B4T4+RAF14i62YrDkA+SUDRSjr6cZHQEzCe
D4msUsRzaL6QkHzCRc/wEKpz+qLXAql4gZR7derxVcxplMo425UDSIVts6g24pTcP0VK80m2lmqw
fKgDWDk5AoeYU6+sipShddNM0rk17c+9l7EKz0uDMrJyIQLJqarB+ZezgALjQuRniOoR0b0XLlNL
DLFfU1/pePAigtq4XrvdsVw8s/2b+A0BzeIYr3RL3m4+DGhEWoFXtGXqGDwpG02EOFxCHDnhe6yd
ppOTlJf9hSXicpZ8ct2Yy6Ra+izQuGYR3qEq2AOll/36cUzt80mgRZCnmMjGlXxSDaofgDTGoRX+
/QvBg6LKJ2pDsaHjgGTBHGNl3fS/LMb2GiyJXO1J2KuuK9b/Ecz2BulCHyVg2rQ3DrqnZi1fuLHY
ltbU+MzL0nMM+vKB/aEf1uptBiLqSJ6/N+8B+l7JolK9TJcH8jAa+wHIb1SWT27RBzUvtO2Y5qfk
jxC5vlYbN5OqLQuFhfTiIKELVXx7qzZMdX3zC5hWHWBLMuguFosJVHvjKSoWiC8IXN5OJPeb3pon
1V1KaDTNdSnpoBXHPtGKTm8sF1VAXa12RTdn4nYCLtMHd1QjEJ+56jXAOJfAU86u/6c8wq6PbQ5B
V4mLRc7nIaz6EF3Yi03LBe/0HcNa/284d20Iyq0ggujW8sbeA0SDuF+PTl8/cqZlJpntBS5+6jfi
b8BgM1EtoUe9hi056YyDAHeJVFPzcCq4n6zSn8y6QytCz9KTNyS0mX6QJNjRfeZ/Z47wkiIL+F0g
2J+ngGqil1s9eD+Tur2ceyVYjpHLU3jxRfvZi0mrXQVxEgezmA/lZgJuKi1PtYauOygsBR4bR0Nr
xA+gsHW/oEeNiYu8mjXAzx8lHvGq8QGvv+iSpY9hyh8Gaw9wRfFiJumqWwlD7RneK0YAHKT1MExC
hGcwSMjW2/JYjPN+l/k1oAw9AyqJHte8Mvgq0+6EtyJg5OxcaRdEmw4D3QRKXvh6f9h9HskavVSi
cP6/KPR921revtvIPZAB7oVuE/ho9HfLJ45yX6UpWUCZAYct2iIEYX8KR6xoaUcA5b6if5Cj521I
sXDbvd9j2dbP1Nk96WkFOOMWwFVVcnHxg+gjwO4vwQ50XDhRdcqT7RImOOFqOhZnxwuXYPZZS84p
FUOU7YJzQnnH9DR5kTRrtP9jM33It5jlF/dJZ+iySZHAIOsMgRUnBFLBD2Rt7+xGUGzbaH807Lk0
4hi7mDM4IxDzEiNy7WUakfusdHnZrRQtFCHx21CnQ9gvbw+MrlagXsFI4MnYE8crcbbADLpSeMgv
aSddAGVURVc1sbFRFtHyMqn+eCKH/JiNCNYCEjBlE+gCYJ39qX+2BDl7RFs3n7Tq5aElTdZCSDTG
jjfvVLpmYoIhIuXHeppkvFjOoxhQDqRrXZjW+eFofyQqoOI87qWBd5q5HCkGS31uo+4+iuuNVsMi
ldLneobStox3MxZlh/2uDkRgpTlRHKLsQ8Ku2v2+2Vm9ISEeoNM6q34J9wRGVa7CIzyqh/nYMeyR
egAs4SEg5gQIZ7ZLwvmnn37956liUfE6uNc9Cq4ews1szA/vWEmC3dt01Rps+de/G7cWQfJ9hKTA
DtQHU0US4FApXOowrLzZQGcnTtJpRIkEdAvYt9Y52HzYg/K0i203IMl/CCRVJNT9YX3vfe1NIpOY
Ah7nS2OZjm/NV8IX+nQcxJ8hRJdj8TgGy5v7Y4Wlwdgo6N0OXCkrkjvtLqHpjKVIIlHYUo5seIQ0
cVfF5lKPW25xwa+EXxxJnckufp7JvfVQ+hX133pCB+0SW9d76ArwSXSAOgtCIC39DNBp0iLVPaCH
DoyCKxIfkum6GfKwTwDw3flEl3FxPHqpFBKGr7rHB+ulIm3hnr/rGKvM0ffk3U+J7JRcFSm2iNrq
oZrVzK6qWWhFdgbCtGsKumogcqQK5olM/ImgqO0RIb9tPxtnAE9L3uutGysGt2V7+Gz83kIIY6SF
F4nSyaIK3JxAb0TBjNwmUSIoevIUg+QRJNlwCB1T5eeYLXevjTn1XXpETY9n/91/WOewwhnL3iuC
T5pZEwjXUi72CENNaUo6m1ae2cM5sRjM9oIntnzT99lIfFF/PleA1BgbN2e2PGATobmyCbR/wP+K
nhMPi4lWAomQiOp2+fntFqeItENd+xN7yW/hnxjEPR0O6gpXNngrkbKOth7irg0HqsEe/GSxrExY
ojscGyat3iK2fUMZwBxVUtsj7QUqLIJyHvlildZsjaNA+KV3L4mq1Yb0juM9M29LQwr54oewag2c
3Lzwjp4Rid0+Rlv30zpVyhQ2kUiiVjUWOlmzT1b8KAEoI7G0U9rx65Zd+LRxxydw/U5Dztf6/HgI
1gpzdLgi73GifgSl1S9eSjy5ZjmI6DUTOKQtMfhU7fThR05bOyy7j+eoxN+0BoORlWuEtFkN8M5d
dmQUPFlkF4A1Ylh5jCC5Z2JyTpdKB1tjQi3l5sO1CqYRmO4//iUxTeiO0xF1bhiB1Pauw7wNj8SB
/JsucRr7fapzM4WcIl3ncWUi/ARNz0OJ7VvPqwhxsYBNIi67iJpmQXnP551TYBiWs4M5s5ZMrIY5
eKtmt4VzECcirAxLDU4Sn3inH7xOWRl7BzrYMj2289RdMPK+50AgHI1+tjBFeWTfaFcXi6bLXt8t
9/2gml7yUiSTT3zmP53xBKpFaTFSZrJi6SOKkCPY/Xe69+iLQ0oqevBexZ/BoY7YLLSyBNJ4w6k4
9BbJEU+isylPh2lNT0IRh7I5fu0EZe6ANsMLFR9AEPXZdrWZJB7oQoPU3Udhtx/IIi3E8laQkpQQ
iA1thI3rdXdAHzYmxWvVFHTZ4xeTtpOiPElucsXHl71Noam5xlsRzD0HERSmvwpwHx0RV0UIutaa
5b4DecmliRXdOSovZBOGmekom89cEsaNtOcdYEOpvNhpTzQUESz1g7Zyah+2BVwMo1LMLZbV8sEc
SCB5UQeo2BozZijpdl3hSRs/ryGerd3urYB47QaIKxGA7Q3s28BgFNHZa0smNgmsq5XxYcEOE2wg
tlGaXVaSDoo/+DCLRSCXm/ps1NCIIA7JheX2mvqCZbnmleUcaxdCQSFtHgItX8Jjs4Mqbvysy//2
MTUs7XXGuJTlA1z3ESZFFK8aO1vIiHQPlF4zMzoMgGQvbp0NCYnaWL2NGw0IjT164UbvvnvFIRTr
RdAuVIYzZ8wpH8NZaUJmkz9ak84XrGhgEMqupwdAbnd2bWRG8t9GTGsOXP/Biw4jQ29ifJbBdPz0
wufzewIx4svYS4Q4lKC0vXH27CwExCAmVZ5Mnts7kLuy9xQZqlbtonv6msbYJw61pPaKDg6Nt8/+
W+2TK5V254cIffGojoUwdDqlpcHzZ6H85CEBjahX40rzHrBUBHjHPG0jpThROH6gWWUFmy11dKPm
wfO7PLHNPlYcNA4Pt8J4zg0X2AuFDbnLVynRjkOEGZN95+chT8T4aAE8vslWB7n517VMqNfK2gaG
NhD+IiuoMf4OH2mkvtxWjTR6Im6+x8VYnsEfv3KAoxL+D9sXLgrKze/R6LIbzFmZqEdF1GuHRDvW
gJsylKM2Ugj9DEEz6Zn8WY/SMlIHezTgmyueTvmuh+4wciFmb/b/XqQ+TSfhROLr9FJrx+OHoJPO
RkWk9tZLmZgxSlzhMtjBw2nejqlyYNjdBc1UVGVxjJqCZBnvH5KlVsaB4WohMyoOBYo3ov7CjaHg
iERlff0ar1Q/9uemsVPEXg15bhAbmxPfDZgYlp9raNUpWPD882NccYRKQDx0raldPWYkFrGEgZLO
bNfYz+KAcGz7BwXVqbhokSm19llV+Z0fRE46Y9T8q8x6kQJTqlOz81oG7GKr2A4yTC2Y0MiIVFOU
q6TAUOjW1Kl62F2iIpL+7+DRepCeqen4Kevdn9ZXzsuBehqkRFasPmtFIzpMfZg8RZxtYhVJ/uty
EPWe1CsdwsvOIHeIe+RPTR2+97fE8SpEtzJsMse88dO6qicVBDiCMvdQtl2I/VDdWaQTzkcuZ2sw
rfQa3B3DkW9H1FeUI74XEB+R6WX45Jij/nrFNr14stnqZMxhN6vFZXEwd5qSzeyUtyZ78wqqPn0H
Q0dNtqWjp+0njQ9WzM+i/bEbmswmI4DsnUltCpZBWqyUJLJoMELPkxn85nFBaBgyi2SGyRoy1eMs
7qiBQAVpEDj5GMs4nxlJCt7SNKFV+6z7cuD0k7JMYlMnF4BLxyum1pVb+PTzkjxDcMTi6OE0MYgU
xYu38nPIEetKdh2tQzd/va3mq3GFypLAGxbz2yFFA2adDqQvDDxhZyqpYLEeHuNKDr9EORHcJoxY
K3djKqu2oKfBZQ1c104Kb3v7bLrNFgAbOH27cpYkcEsMLJqoMdRhiZ66nbFXzB6SzoODxWybLrJw
bXQ9uL7788LIQKsW14bcDmcSoqD+82pXutzHdG843inkGlUlREblZuCifnGI49XdFgHIgKUrZ45a
hhL6oUpKB08Z/og+uNsGCYyIzUlNU5aD4lDGpry12Y88+GKuJgLMyLSgdyyT/R9D5QzeI15yXwpD
VekGaRy4Cbi/BPzmdgPlepJHvYej5Lh9t6mmjhgZk0zZok13TmivM7jpJYoHGRNZRAidssXxS0lo
kvupYM3Jan/TCXaCAy/nHORqvZr+Xh1FVY/jejb4agCdl/QLBlKq5sUQ0ZY7h3gEme8sO0zK81pk
bfZ44Z+/BEiwSN4rM+73d+0ToLcf0ayvJkjndhAOp3LIE/Xsy06nPNLpwZCTI7puyDx4plOkWP//
8VOlN/+edBozJONFEY3aYua7pOx/0DaG869/7oTHCj6OKLS1c24YROJQEXIrI8CUt1v6LDGW5+lr
+qjpCbHhMIBcYDEqmgJRksDPFQXIPIw55SSUfmQDnWmR5NCFFEVR/JC5khCv/Prx4s23NjvRDe2v
pTevd+5SJKV6JR+D4oUTbTfuQXh+0pbqHTs6UcZmLiwsOhAi9Mgv0H8T0am9yNhYCGTH1AJITSv0
/sida+C1Pwx6ZA5hUbu84fAxFsZpIWJ9iQ+Wt3kRrvYU2mS6eKQhGSn7SfwBPZTNB8qzxw26C5V0
LgysPZpKNDkSPqKM5kWLf+kk4yL2n20+oobduE/tn42MFS1QAjFGh6isSw99teu7tsP/F9XI6bQc
LM6bNWutdNYwCJGvP6E++HfCXZmUmjhnxEjRJkH9XmQkXIjr8DMNMi/wurFy3RzBwBdbYtN1TBfE
O0XC2hGTxys0Um8wCu/NomDwgXKRDxQUdwRqnpWhUwoZbRU46gvZ7zxCRWCkll+Mx6ApVyProdvq
NQhvPBgUxJAzmwIbQ05eDzXn35wlzBaYOwuv1OH0mbHJPzXZtvXyqMwxlRuQUIT0/UXiueoubHIA
g4xVIZOUtBstN3g2ShN5Bc8AqDPXpyYdH+cUvRAceC8Tqrh3Xf07Do7zCqJbdLz3B3kZBxWQ2HdH
mPErhf/SEB06ksuXhxOb62qA1H78m2pIkt6uUDvFY60cir75RXnRbVCVYy4AYG6HBWavDCBQxza8
3tyFy5e8s4QBQdeqvZPQojV3bZ9W7GwspY9RvUbGWl2Yt1UFoPv6mbp0ekZFZY3gBHmEqLbjG9AB
/AJZhVMu5DiU9e02/jCbgJTtHj+IWO1TbTb5T6vYb2sMkRxn4IoqC4pGHlPWf8iZd5beBY4273TY
gNU9pnAeB37uXwLYI7vhMMEuKJJsNkC9+Ku2EN7YZ6iJeC98TnYIEZJUle2thhGApStx/ZkrccBr
OlQjGugxGO400KRTFWZNLjpLctlmydu/e4VgC4er4w7rP4axjJzESZOn1q8BcVK6KFgIPyqIh4+O
cOp3BwVdVVWjbZA7SStIdpA8ViLjfZZqAQhrvN6vqlbbTGx8zFodGJEyFjC7dvUeoX3/q2jz2jDB
89mx9Le23K0XLaBdmbkJEbhEIDNGorxHGQnufhE6r7bBWprKqssji8aGfuLl9KbxtCWGz4Ntymuj
L9NyEB+ZgrCCy67Jeinu+yxl6JOZ5bT7DXeDSiMhpnQtK5isolaNG/9id2J3B8BCsEFtkgUcmTu6
nain3L0XmPx3DSXbh47SqLodPUSyE+oNnhwjzxVkL8J5Hc4U/1Fh1Qs+IAch3XqBGAr6rby4aNCg
U7XN3RGQkn79fIS105ozgUv44h7abdho8NR8B0SOJKuEOw7zhBZ8ESAhYEfXq5xl3VbKgU4yEqll
kQs4BkZyOlcLeDy0WOaFiw6Qi6fdkElvfCrmuOLuhx3//4hyH//10qYjlLoZLbjCaV7wXHQDo0Xj
Okl+nLnDmrdVqPaihO4UCLDg17FSx5BjtzWCG/8fgoNWreoceaKQ4LtjW+iLkdH8B1vt+ZK/yCrc
zVvmWLCUY/4yu+bHl3EEKVKMYZmQUt8o19L10s35qgPGtLeDkWiTuEy5QYY9Y0TpGcERivFFSqCi
+jnybG27l0pY35QbX2ZglP9F2h44pVlN7V4SS9pIBS3tNCiZ1e/Xr7xaahwN/C09yr+dI6O66Ioe
Tp8IiJtJlZvjUS8+IcGayDb7nYoZsQIW5xtkU07NxTMUo5wM0vl4Qfz4j/TVoU1lr9+mH5LM1NZs
3cQ2oFWuV6EcoCjpeXtEh/PhnqrsSNkdD1vo8hMC8P/sHFob7z/i6qUZ3DyJMxtQPyiglyLKnX9e
F4kG5bV71dlWGeI0Mg27FgDqeWea0YkiixQKbmkWIysrV7ZBgl4857jHkDf5fJJ1CXmIodVrhYfb
XigEFe4KdL43I+A276R6vdAZe7FXhIe9m9bdKrpLMGbf/dwiJaeCBGKfz77zB/AcwHY+ck7gaHrz
CS7zGRp45Ku5gPdCYVMv9rM/Fitc9jYNThxFjugd+AtbScg09IpeQjY5I8tIy8cKs1L99k4bBejv
UqshX6XDdY+0I00PeBjdCB18wnJYMuDYG1LHU4x9dv/rEaZY8otLGqW+hkI1W+XyPubBrYSFtEFF
bBPYhr6GPGBzB5m5A4Syygl6W4S1549tWGYvRzV5svqBBy6k9t4eQVlk4rL4KSYfLXNKizOyX0tv
jXU2aXzeXld1ndpMWl9QRiFsG2Qe6jp8jvieljctVFHWHjVsI2eLOfXEIRDKIVTXp5l91mpJ/w60
4LRQ+QiHXjanE9XiY9YVu9rqAXY32h3MSkGw2SlD/uROv+YU0NdXA1xfb6zQ+WnXfYA/sSWLkwzn
6JL4Kkembxv1oIWSANAh9407vahDbKkM3Jx9jDgWf+wmvvcw7wdcw4L5gmx0kO20A7fgsorDsP6W
M0PGWT9tfKxG+yDNquu3v7Ky+U/I2cnLxRnEINp7VNHfec+d4bp/JF7lGEuh6aU2B48vBn1CzFnL
0regr6/c1XuK/tH+AYeBf9mdxT4ZPCygznlg5EPP26H95nIQ/jSLKCxZSddth5CxpPnhC8TPqaWy
uayRi/pnVWW0ztQMzVxb6YUWsHIO+4s+37xWw0eG2XOVOlyAM62FvYXofiYFthW8FfcBxEo8ca1A
vIL5qwMiEe/LdwJdkF87Zwm9sQgWYvngTBb+K6iwjhP8gDwEbu6/neo5yephX5mU9tz4P+8uF1my
9lvR6A2gqgkeoUGe7tAu5XcdeKHW9Sa+MnVWIg4kCSVFY0IDWm2iQOQ4MGje95N5TpMbcLULs26v
nGRbLtE+982TtqV+WGd2YwYMg13zubzpGvcF3W+OOANHyd1I41xG1WPlH/ta2q70ZID5BRiqkGgV
G0OrOme2OFsCOZJ+lc8xMoCRHzb4I0fMtqTfK0BHGnqa0eqzfQUj4Jd+Lj1Kfe/+UfB8JpNSRtuS
PdhONiyeYuWhii05Z71sYdQpLUcKwVNfWJXAO/NhnDnJzjwLWzGAooX8UAfhBDLEOhXSx+zPajrO
prCgXXY2s4NeTupH+TzluhselELuq5pBlAlEWPUNAjeatZl60fbdqYN/Vtnftw3t3YwKB6DW/rom
aZdhINe3OVtA4K78JrsskkE5kVFEbq6XyWq4cEZxYMxXF45RkHI2TfngB3ELMtOdVxjCw+Uyrrad
Hm+dG4QYDMB/NDECr+o171+7zuhyI4cf5JWwV0xHSOVy9jBBrs7yz9oElSU4nCqmIfB4SEDTWRTu
jOe+HG9Dwo35y8wyQ6NKOE+6APDPUulTOcQS6gGDZExp33G79Q0H5blzrDODekiJpEUEKVwJtO/P
C30uO51okVZfSjMJ5rICR1Q8tDM97chWncAkTW06+P1hHPb+oVOBQdfi0sVOI6wnveOz4++gJCs9
qtGRg6NJkApDi0Nv0ruDoqNWqgozBxDvXPvqtlTXKZfVjKX8bSnsaY8D+xXK5RMvmjdfFhyXJebz
6ecvJondGafAugeb03et2tOApyP/JMcS7Yp2O5PXNkix5vHm99rm0Ish3QHI3FjLG8ZOY6TS7O/V
K39jCt4UQVDD5xbcQk9jn14wguFh32edzUsSbtLYVdzrgwdRxdrjr0pAhtsIcHE+M1v2WKP7pWZT
GCiloktIMd6c+/8Vketub2JMTf02Enyrj7v2epAyPc15+DWvIskN+ROJ/W10l5fsZnr3O5YHHBjR
pYmMImNJaFIyccxFFOWeKSd1QYDO7lk9c5VGOWY7Pr+IkjkWJ12a0dVRUnA42zg40Ql49s/1wUy/
bG5YR7D1EmbaAG1RAMosn61LgJdgXDZp9Unrt3X7Q/ys7sP21AXx9UH0qvzNECpWU/t4rtnGPMvj
r0Jeat4Hni7bKVYZQ7Q81nTxvfNbL1+zELvU55symIofnvjtvlTlk/tiP1mSV+EcLu3RgbwaVJBH
zes9VCjw6HtK4NDDkOssuHcChyW3BpsS+sAyvGA1vCz4J9UktzKhzLUPyNbWZj1ZRNZdRF0UauZ7
d8tLAMlQwEI7jl7DBCRVRTSuVyQYpZXAz/7pTFyAh8Noi3B4uQ32mB9Sgdug3A1xe+p6/idgCfGV
2MV4lKHa7GvdTVylF+juWvZ2bNTGigMtuMuAJ5DSCn1IkciAvoHJXgs426jVuptVXNx7mFu4pDjP
nH4xzUAqElFWmXdsX0PhTcZyFRg4V/3WtjNG88FMrUHlYWdCzhUsCSOWo/oft2mwVdXaiBZMSTGw
WXceFDvKs0jIbd+ke0cYUJsif3hJeBYHNIM1MvPCbC+pqjE9efXMxKousCrRYf0e8CK1ucZ0FV4l
WPYFkpr0KFi0EiZnNR9PdaZ0QvdGBVaX1oCPmIqCBSqzgzn4qYgIQtiQzlFyhMYm45miF02xj7bJ
9gANzNQUqgdWmeKdB37hQkQ55NmQxPFDlHtX7YDC/iDmMwNvs0f7D5C3ScS8zKYkHvh+qNhGGbXC
BZwmPE9wgoxNDl3f/uaaG/Mlf2bppe6OMeJHu0iKYn+qK+iVG+HRazLRLBLL83OFk9zY68G4wg+1
2yBeXTyQHMmAixefJjr/qBl7Arwmgj6tGUeUICvcaLvpJShSgY4gKYxwtUhE/A5j/P5FfeJFOIEl
aJYvlege9HrYFKLaIpxoIcbJShZQisu/UEfdIqyVVK7fIiUOPKT24hVo8RJWTdczSPpA1X7siOQj
loOdOUkJvX5/Jb3tX52a+yyG74VkNfY6P4uOKnfm/fLHCa3ljapghjQn4vP7r9g5QAHs+yvlUd81
7zdJbSQp8LjaCKzTa8hEscXGB0Jthb6PGmjFqWpvltZ+Op5rLJ2A5dgm7OQSEf142UgjRUqvSW8q
GsXFdvEIyh9z4ocl+PzDLVSLNwraa+S/SwuVi0PrBTUeVked+l2hmMmsdEB2tvl9p9c0h+++uqXp
T8s2cDvWt2VlG6PS5OSzC4UPGDIR2G76Z+1WmxmAVOinannO5akMdzqucVTy9M5Ey7QVH5r3Kc4/
zr/7Dc/tYESb28fZ46Mp9v0W68H7KFVV05WDRFsrsJYrk0ebL1T8aKSANIK+QUSpnX4AAPes51az
lzs0qwFyQnKPujhY7bFjPQSzEp9KdNIIOpmYcauRH37079e1FiQNRHqy6l+LRhHCB3+DtLM8jqmR
3EB71l6Psvuc6yh+oZZYWwoejYJSNr5Y7SjtOxz9xdRA22of5qJ4OhNpgh8DD7T7NChh0r/znQql
QPVsiU6wMQwHABmDV5xIf8xHgf9w48HX4PiFxxxDZ8nGeycGXdhSJe9HyokkSILeUAiRcScPVmxx
Z4bF5Ue7i3/VW3AdPiS0OFWVn6/bK0vtCDladje0Vk8GkmUZ1H9Al0YiGgyx7Ss06fDjqMPtgm2D
vtBs9mGMhqjcMYJ2masrvoGMWSUJZ2ytkna0HTFV92EcpgBFqmruzv7LqJqFjZC7UWoYktDwsgtP
Tc2bQiSRY5u8ra9ezwTg8aIZPeEvvNOPjDCo0uY1xeFr6CYA2HmDcfg4EVhwpshIVvXLGqq/vBVC
V21o0Ru4aFJtgb+LpylBDtl8kRg54fDqZL9V5lrSSo3by9isBe4iA9VjuDFMCjkntdWzzJMTdata
bnJ+TTB/PuL+Fw7K2TKK2U760LZgats/eo2i4SAuJ9wfhN0yWJBdlS+4peWTC+o3OQYb1pNFVOOH
cffhNFNoXK6E87PE8Bnf7z5GT4/De3ksnTnUIBX4z+wL8ZIx5Z3PKm9ZwNfgKGzBhw20nhvF+Gi2
QbdQ5d8Pb++Szvk8VqjsT2hR2HbTX7KpITROEWao7yHv75mJTxQvP1h+u5UtVWQX3G0MNNUeSlrJ
6CBNuF6bfqE4UUKAD8lrr6GDIb7f3WdtQex0+u3TkzHLI3UemxJa9I8cs7WHNM0QPfC3D0W4/Xy+
SNNKTu43C6jcKVp8TKWCIlVFfMVgKqdPHm32Vl9USMre/BqL2+zPstfKyDaKBQlDj4X7A++Sc06M
LjhXhN0PwTvYWLghtRoB1TDesQJIQAQzeZhpS4RHRXzwIzu7+cn1hgo7RXUY70iTFWtEALiGnDG2
d6Axv9FGNG8gPKdIuvMWTAF8iGPUUxtR6FJqe+lAilhZ0+aerCB0FR5aGZg/YgrLB4AY0J9wwI2X
sh3CyIpCdgmoHkxqdM23Bh5pyhb3Kd5Qv0cAaMWRplPnIsazOWd4j8YTKr1ysErWX+80synVSdJC
6SxWAON0OvRKfYw4dz/+HRryqJJZrm4FZnBcqtqMg4lGSOGWnS8wIikOSQ2RTsELJzsuZBJzCXBk
BovL+jeN/qBBfFgaZFSMoi2I3GSxOCDDdShqeAZQ2pzfxKLh4GyH5Kg9G0DKGxazttNPDrl+59bX
6rN4ebsGf7fs6i6XcTJU7eZUPbLJTEGNRnW2mCKoEAMXtCbHDp9IefjKxudO5f8af8x+/uzh5CD+
QMQc5Ku3bdJRPIIyCPMvWsOTHhspfX7IeqEmh0y+xMBLgnwe5K6Rl3f6kx5YFRC+EGNTC7BV8owZ
SbohTgqiw586C56hJtNkEOGpHx6o7cALuOZYKpOhjZCDl/2H3eT5JT6z/Fa4LBeypt6LfqJ/izS6
TB91sFdqwNDgs7ZM5PxExzURAg4wZoURoRbM2laqutMlM7xITYuCCI8s3wCw2X9lLDYYaTHa+9p2
9y1PRUpP5qWEjJ9jI9t5mQHegDGXGKesfi24d+HBgjE4eDxgGOOaAJggX3fxoe8YT8Ht1PouGVdA
uFiJ41siF7aZmmzJhA0JTPCsIPoFwQvtl/5bWc0IrmZkD1WfGegJowIiqwLf/t2WAbEx/0hyZmB/
Kk+yRiKp0ROG6cZQZ6P6sDNd3GMlVn051eJKodb2yXA1yA42zzuVT5u+rAvfjiZCciIL4cK7HPt/
8+7OKSGOQPMSzPQdDz24S89v5iO3eW4WqiirSHPV9wUdFKmYhS9TWjZ7qxQK1BfnNsVzVq/M9XK8
UVwBgYPlkihV3seTzlqQsIsYQghZACp+c1UHihd1TQDXmPm2wbGLAxsR9eikRxSkEZ/tmOlNgriC
XZJQHW3DjD6VF3GYpaDM1LVoe1g5LmA6gNOtEjQSwaH/u2vbhXhj9f8PtBZM1w7CmCgXJIreA2AZ
NRINg7uSTCqM/e+2098LkqN4ze6M/o0Kv2VwANAVXEAMwIAPtcz13YnxU4FEmWRLrPIVC0SMvse/
kK3jFE2VxBmBpvOYGh+XYEfUNzy3PHdi4k6dsiT/vIZTSstA08lP/spBy99673lomOJ204bFva21
iVRarpgf7+j8kS3Fd2RJIWgnfQdr3FAZw+bYCQnDd+P4CgHbUPdixtGKU06AK44P6Reto1bg0tnm
iTjcWVBuRRlTLDvmMhDVXJyIYvDO2pHVVG/PE8Lmri4FIXAwLRhaFWfa9K45Xj8SOVSNlkdlc6Uf
5gGZWaYjyKXDxsraKgahZVzEyVlF6Ck/JW1g5L4HfIKW5rU67P44ZLvI8T52mxICCF29ez1VEX9s
FO6Gv+poDl/hUObKMYALWT/uh4hEi5fgt2sPIY24toVBRZOAj0qjji+/Nt6iS/1QAJ7R8kKp3r0F
yX4E8DxPl+SLdJ6sU6TTuR4NHFK10qsgR4O4ZJ9XNdYtVJIWDfH+eiMjFBAo6hS4o1YNTP5RLbF4
YMumeIV5Ud+7IpWlR91JXQk63EROAnpW8o7FvG7dLHEyuGp4XuKFVkB30hbB016Q5cyCP5UzmSKI
XStiz1v7MlLibpNUpulqdELCtTGo4PiS/MAc4eKBw8v47U5B6Uyce8FN9Uaf8GrEDr9Rb6yNixmE
YqUgyYVKYqMGJg4pRZRSeD47+e21K6bSUF3BJOa4Ohe8f/p5IXV9oXE9/h8Vu5lNUleaNSbXcAhi
iGVTrE5Xlr4Y1dv+6CvPs839AiaKOHHyopcxuCaOCrLgGZA9TF1kZq0BeihrjgkpPVQxDGF7FevD
391paQeZ2s9WUMg2LU19Q1qkYVzLXNlDSLFkM8KkTuP+XLYF8SrvlxyIpFM/Rt1gGWoVMU882A7/
hkVXbKQyM+AgS2Yu1h3Kup3aWHEvVML0Y347t7g6l5OI5wR+I1oHUb9oiZwi/JyMSByetdkxhDjs
2uKmckHHWbaBYCzSVjXH+ZGnq2U8MIN5/TW4bJWQekz6cbrMQgWFI2da1raBcw/M0F4GSTxtY2Re
AzZwMuu36uIZFAkCIwL68NdGwF9XueAjqEZ7eL145QLAPJn2Oehs+KAR2xU9SQZYFhzX6+bOCXLo
8adke39kv0T3t+yLTFtjMm+ywAVoB8otfOMZaBzWEdl3meBn4Zw3oueX3iAmAY2ZHxu8UMkte0/7
6mYnR4BQxPGbHhSoj1hC4fjvSPiY2YIApOTBqtM+ueYvKPoMqUHx5YFfr/a59v77pLjoEW4fkMXr
3Rf1JmYOdaCUua7CvHOk9u6xt4DBr1ejXuaWloCpT4Zsa7xl1dW5+Ks4dfpxoP5zEjhWFnr1H2yX
5xB0+szGTZ05jik7uvsZJhewyqzCd29n/ILOyLMJLZHV6f51ohkEF74BPHse9IOydpBHCPIptDCX
IwEBZlq1sMgVi6pM0pxtVuWZlQ4/Z1K37/C/WSsWTPbTa4cTiG8Wf5yOQfNmdy0cWpKIfC9ESsTu
kZQTcHNs1SA5KpeTesHDdpoKKagJS91L5KpEVnVjiBDPw7fK4ZMndzyq7Y7Dwa3FX5S/YSMpkdM0
JY8+GSrvWi2VvgZ6Qr3QaTQvbFfMO09F0S14GkiHBGlFyrldhqKoft3F3RPAAfVxpy+lqGuyiyqU
bPI919j5sRCwxAPp0zAY/8f2Z5ZYQjzW3kbXT8xA1wSPvcFjbUN++kQFQncx24ST9xcjfetiPnnG
q4TzSqVx7i42/WDhjcP5N84RW0uBShxwogya6ICPBjWh86q48T8SsDL4MOnJLIA58I36/zGNLxnC
5i0U8KQPwSOZYJJI2ooLj4xjtyZuTDsTrtq2MxbjO8OVuG/KTVb2Qb8qMW9doFP8B3icfTjRn8sz
y6zx3DR3D9Fuj5lGK9AwYKV8v1AlsVY59Is29d1it4TJ8BT4CeBBeKIEtTNgb91FGjbI7zuSRiRL
YYBmyptp2ZdIyDwKuCQybB7r4DrSnaHw0AMxx1yCV2BK7kx68QCDl0klctbo0WhwtPWgGlxzG6hJ
Z7H4LgYJYPKaouWVe/Fa11izCeFuIMxgh0xbtagDqHlpRbpIPQsY6nJ6yCSsueGHEYH07akLF4gR
Bw94RT+JEH4jQTCFN9w1TbjSTUgOJ8VzYrfE4gPgfes7Mvoa6h3sPJkTLAEKDial/Zh41wsLSW5R
9ZEfXeMG/JoGD0zFYcoz2FEc/51F4KuD+bWXX5lAIidsq92Bqr3LhpanlcDx69m+7FQaSw6H9Q15
JjJ0kfqxrfYK0EgWQ1/oKZ0kNGmzp8UmHOdAz8i1cFuGx42xXMyAA1lXY/CZbt7f4fTMjEMdPmbX
tSqa17RBubKqS63ZA4IA0UXE1JlgwtZJGRdX2tkdBRh1FxohqzHXFMDq6OuCQgN3u/0SOxOX2a7V
MxbkgbvfHNBBeFnG3UgUFR+ttmeRbwr8yYCAd0MDbsIs0E1xGhIOWC3oWqLQk+V1/Y0GpoTFaCLX
iOBK0YxJS2CROcy5+rhSiXwElpynpbZgYymzTpImzRaJpgg4d0tAApxaJFYKfMQ4jKNZXZ9wZb9j
CEWplNwVZFMkX/JwB+tVH1gU1Z3IOhMcL4F7TY2WYPxlLniD3tdRSksJTXX7xlGIrvOUTJRI6v6u
T+UhBOGBzGYMuYAz4JKV8tZtP1Zaw3XTguodklKUkBP/ccucCUI1N0e64TB6S5N2lceQtC3KPevB
1KeDKvJLdwjR15eo6jrUk0oHY03fslte61KyfmRHgjFzFkb0t3C6Su5leqrSG5v3ayTxX09PQERy
pklbo2ibb+bOcn+1UDtCNaQZrnuIvNRX8mas7n2W/oEzSFdZGtnzsRGNwGrOJYbbhyy+GzZTqF9I
+yFOJ9ZK8L1UAfte1JtkQT2UzykXKuRhiZ2cP6hoChIk8LUfz8GTVv+ThXSSpwHMjXnD/40HDR9s
vhU+abAXJRNFGEo9tbfk9mmK+aScmU2onrEIkTD9j5n77H6+pnPS2ePEdWaxpu8YeQcKPH+OL2y7
cMo+6gK77MtBs7dzljT94xew9Ey8PIoZhCSz7ZCx4bxMjCPCbEDkyq/rLWxhxV7pOBmwpzoHYUac
7fTAxRPlxX4F/4wu2CM6f+Wv/joFa1vPfUjhdpdpaukBmxtg85cnxZdYxats1NYeCskdlmKvi9jK
KXkwKLNnuBiAYe7hGT3BJm78vc1NFTJo7FwHq9soz7xh0DRJTH8SFwjN6n2uxrooPcFf0VKSD+Vv
9aRAuuIq/SULrdh5XpNrlQNDpMPzVgVf3yM5jrYoUIZNmOVUqZQCnjS++/OPTC8F90m9HUSUYZ+Y
Ivdzu50Bjw4oknOXr/V7h2iu6SmG8B8lFWayR/ie4VkoESSQLgziwr1/i3ifFSztxDqnCLeUvpnM
GDUya1A1KDbfRCYqGHKV6bhmLkQF+ptWYcJxxUN2/BhHXYAfURp5kh6O1AWTDK+7zMKJ7V6dHUbd
gS3a7s9Sk0sPdcJnWQYHGt3Tpjt599/9/2U8i5Ezi4NzTgS2kKLPtHa5pIDUe/Jk93j5jTUjSkYc
d11Iq2mZOvljoTGwk7+e2UWo8wM7j7mlBVpq19TfP+JD31dabXCC+YH+/ftdIoA4dnvOVzDpQevf
2lSDUzf+HjJOjBL/0Pr1w3iu9RnDpka91ECP3BHGpG5s1P5XtEZKPAGN+W+cCHm1M5X5p/B/K9gB
2WPHotbKmYt71+NErrnNIF6I26nU5G5FSwM8vdWZANMMltrmSSKfvlYCfIDZAfvFya8IXtE0dyC3
8TrplPn3FKPNfbhCN01M5nIoMzAp9lQvl0n4Hgva52wQtJZAMuVJZFipcHPxGoK49F/TgTEi/tP3
rlDbEbdexg5bXEuqoVEriyzaWQnfIY7u64cXxu9y9POxD+Y4cf1lawd5pb9Y9pjTbR/ZvE9Zhvwl
WoY8XlLd3eWqVm/iE3NMTJFLJb+7hMBJRbPfzdHmHfUXOI2LaZX9J1o4eqPOndrcFQ+8IxWXJEDb
8M+5TBN9+OJZWBNDBxsrv9xl0C6s70l8V4rQBhPUUwYfEnBApxYz5iDQKVWdQWyTPh0uSVQM7521
RRfAcvSsMwxsfBQUZCEb0+RK3NTj5yKVwl43vo+wY/j/+cfg6F9217/UO3LQmghyM0OybHsRxlpI
YtpyqG55TZKqrGIVN61a1it26w6jaZBo4slyMz987Mvg3d5qgdFxEqRKs7P5JVVjUFcJtrJMBdTK
rBtNmFPKneltuD5K2ydPC1gIHa4piYvQ1ZRaQXwu53RHA0etJbl8YiFwnRbnIFsPeRo/UfbZDiXN
bZmV45ZqG10szTBViMupRQufZpujcoo8HoKnjpfMHQpQbCpFR5eRmEPjNIpmyFvI3WUuPkBGnZ1s
BpoE8Lr+sSCx0VXv6kvtPdg/gTw8JxodL6vQauIOhqQlQ1tBYYiqvw/dBUBl7W41KeNce3eP47tj
DhPRSwnGwRzbS8SYGhGA2BNI9TSjhVQOECnUf6AIGfTWup5MXdHw0siNAwY1Z4zArMpXnbEpCVUW
3TpDkIez9JrOqQ9O0VMJHJAShvHRzPVEwXsLp4bjUKGX7xlH5a5BQ9JIdTNvxvqQD1vzF5V0i9Ct
qN6wftsizzCGFvSdinOrRoGXzUt96mGGbOb5UJq5536oywQfp2XfBuc+CUs70EoF7KwLF5c24W/0
ld2uSaQtFRhX0OZ8A7FU9szvTp/jk1tYNB3POzfsBiGyZSqUJPSW/494tOCsqsFSU9TLc6rQ3FGI
60AA+B5xmVv+0icjxaS7DrcLnrBBqjxNTvmxzDhSZEdY/qTOihoF7+O8Ie+rv1ijn+9ekH6B/Qog
H/draIS+NZLesB8F9xUj1PT+BQHWJGbQM7zCjqZ3oxc8Wp1eFgaYYse5MwZ3EAkqvTxbmlLY2EIQ
XJQhJuQ2X+OBThNYFh401mgAGMGhiK+ZZ+iL8xNlCYu9voP3Jz0t2Iqvhqez+iyrEkU6ahNXGMq1
tyI1uU5ajZf4p+vghv7MUtn3IQmB7cG2jA171a6EkHScK61641naWMNZtpeqF/w487al7mT6s9HV
MzvjRnl3adMv5Uq9iTrFdlcBcFd7p06/r9EwXQ6tWvLy8F4rGxDmn3OdaHizFhMDQ2BDe/Y3uSAU
j1j1eOA+Z1Ah/dmDJ8pQFHVVGbPIN4vMATTe/7qe5+4E7UOWGceZpq0VmOvA3Bjz0D1/TmlxQalX
/ITqFZy7GbsFt3yr+EzqMNcRngprN2oP02rqm4tmm5AP8CjkVDXximXLDdRTN4A+fhMt6gbk+0Ds
caB3Wchmga4VrTUfOkEVx/6TYvXEvuHvxqMREzhF9fD6mVHbebBq7y+hnYYREMFsTf1zZdN5YIyt
KDqQAqQvryR+tgXkt59ff4IqLOViJExAuMi9Ry6Yuv8LBKXcWeqi6tEASCxYJuH8WaayrN0Dly4B
OyJ6KbGzrNUvPwjUO7jocsaKQsXlzGq7l/D2ZFZk2Fk4fVAk5uM4IDThpByW1eVhjwuwfuGH9y2e
d1p0hbLJbdFBnteuGnJr5d/PpL2DW7Ix/rWlwsZ9bDaYcLw/UEGkS/c06Nlhj1AlzoxEeZTqVvbz
iYXb9O/77qIWrdP3oXoNuvu6vhojaPrAL/LF3OfFHz51UmAvv7t9rGGi3B94+NVoXqTogZh6Ebun
01mK1YRffti8R2L9ybJcu/56LGQT4TvQ2UDRYocWbMIuIQ97iPpGHUitHsfBahOESdr8ogUnBtGp
NHRB3LBHLzSb3uuFncbrN0iEv1btZzi0PZh6seleSqIeHqvcKlXYxuoM3fuUDW6PtQ1exhUxf9bB
fSk4IoQeil0NVa6TrWm+4rdRRBW6DbLqwmieVTRzjqae3S8Zxirkif1td+OcgkfSCaN6656LhyGW
tJ8CqJW1O6O/kMY31MXNBvQg4uclroz/GrxSfBOtN+8b6tNND36EhhnyDX+c6IT/5wjp7IkPdiu7
sOxopPlJXxdnYbcFdizoV4xEb48TH6BRhr4RvYPDXL78MB5W7VDfRQSweTKerXalN5cHvv4Y5ed0
45qqkugSju+lN4R/XKn8iKR0qB1rh53RClMapv8OmZhMGXe0DL/mwfNQkr9w2rwOGdadBH5k2Pj5
2SFcCTyFi4Xh1TOb2K3zJkO3buVS1/ganyS/BNRd0nKCMdBk98iQUpKnkLLa2fWRuFi4a+kcNdja
rTx/Z6sPrEa8zrjOBU7AUU0v+aovrxEeU+QwYleeObBv91hf4vAn/ZkBnDVKsTlKsoLoz0pjUFgJ
X6O+7W7LLBQtMNlSywhUK4ymOTFilW3/pIbe8bqGxBU3d7jsXnpjX5v3IyrVZQMPsYh17HcFnqee
UoIx1BD68bnGRJzlA/1qSMi2BAPNG/1PcQAJfAvW84/3M9OClrq8830KvKZ+NVE7POLLeO718h2U
Fy0ckgV/+RGO4boaM/2dl7TTrFgAi0vLx2eGLIfcJydSE1IoH/em/jXPXieRE4OhwRJjR5IY+qxD
FIELo08lAyWmspAkpYjRhaCGuvVi34XtgFXN26Qga97pljchkKlJeGFGhdNSBF/QKaLnnd53Uksb
aACtlrI6hVx7l5fhTGiBqr899dnP+5fkyF0LOf/wm7R3T2Ht2SACevDpgdxYAw5+bXiqdQt/+ySD
0nLZ2/mJ2UDn8DSj09EsTTuOIeCaAUHMjxlRWQ8JgpF/NHrt+gpXDbULwxushcOAI9lRd6MjJ1I6
TnwVqhqhTUlhazHfzKxJxiMWy12lIs2TylDZozNj8yuF6RvoNyyYyezyJN99ZThtxZQietVgezUX
al0ODxUzxAQXwPzM1hPhvdeQshd4CYcWcS8c8DKionTBz4aZhnyh+rvUlaW7LHpEWGECySzjELfZ
sZDfCmBK36x7wa920B0m9c86ds1TpLCKcaXDH6s0zIcP2uVnVjlOGT2RSkAjyBN95j64D/6eWk1l
GlB1U/BJUkPiulP7bMFAW2CALKra1h6f7S9QicWt2KTopZMINM1XnFtNruzICUDBZUPG/gEKrHdn
gDh6qP9tlJoPbYQJUpJR2x4mugADDnmHV3SGDd/bB9B/hu6lfdkSsPDi3XzBxL6QkUWcKToP5qHs
T1Japal7LqKQbpGjwBoDwaQiApdJo+jcGxjiGvlLSDRmBZcpbOemnFY7qcoVde9PXTk2QdR23aew
0wXb5IQRLICu+pHhMjQzWpIIJwuZzVSiPXhLPF893SaNv88lNyW4FpFAICzmCQ5f/oKv+bR4NK4K
bJRkCHlcKUwcAq3N06XgOJEfWE2f20Ag5i6BfAAcDh83PnCvShqUuKEy8uLazN+ZK7mVnvWzkeqz
z81mv8DJAiWpYBcTRxO9Z7sdRy/PLa6tgF22M9LUAcCOAunIZBjUcvxyjev5PJIUZyHm1mqz6XVP
wirrfqSk/LfY7aI6joelj97mjdV0LqdpCW6w1r4Z32XsALfb6xCfOTSuP1N6CcOy4Np5U2PGK8Fz
MHgyLpv+yiNth1v0VGfRDC08+Vr675zI2Wz+k4E+hXLV+wmRronwlXiT2olA+PAO/PyyTx0772CH
pj3Pxy09xXiVOdLT5fjEidSMuBRd1YGYym0ZFQRScFxS5KJGv417+tKd8Gtfu2bvQkszZmZjkiuF
MEhSRMQQt/sFxDoPUOQdpuwxd4MJtDWP+giczBIswZbKPHEOk8UO7gvO/Y6tfHeOAMmr+SPPzuXA
BBrj3GxfiI5FPWe4epAh8nSrQhMhwcb0+Q/fQznpssG8ltHfXFYglRWlgwWqV536GbajNg0wVUdY
aEHUCCdfCU9fNem5ujSlE7p0FervldqCPKCdaKhzRxf7mXOKIn1OaMRdogxSl+3uX/8QGWp4hrm4
90btM8ETIFekFQAKIwlPg5kb53kgRHn7RqTgTHvhgzr3d+xeWbu3NMXxTwBTmR+Xt2JHcFxRHI3r
Z8R3WfL0DvqatEn9vZgWAo/UNNJc2LRO32ibEL66OOqieJxxKPhw4TnpHWjzzCK1rRssVwYlYs5N
c020/fJh4bSkEk1AOtQ0K9tCq6csjDrmQ0w1OCSx9Ub6nbIkHI9h86t56VvdqcLgV/XOd5E1CwX7
r2vP2UpH6IJFb39NV1OSk8rO/VelDe5XK21P8QKtrIbh0RIj83/POcZSypp5u27HmNqLVoeO0yWx
SKQXlUm1vNUcoXJo6ByoMWbH9Tx9ZSsr3sq1WaeqYyDABsi6gYt4F/rNh6MBpN+z5b9gL3wdMSEc
3C8+bRZPI97vWGRFsONZm7CGIEVYTi6X1mU5s7ZsC9ZObHyGmVOv3uK+/x6cxWtVza5QOZ1oKWgR
IBxDaP1Uv/gMkI/a6+wIFexRlCMs1VgOM9SyQn7M597XiufjXHjPgA5yVfaAuFw3p29MZtquXpTU
K2mmJmPQ6eh8ebx5oSfEudEuBYuMdGt8xxoEh9h9EKub1am6Sg7LAEp/J5+AWRPqMI1gRvVoPbQc
LGWyEGkCP3zMS0eWaFqIqDJVw1PWwOfUE8kfvGYHb2/ajTA9vF35BZ2HUxkpzXO93pnkcBChwSos
UNkZCO4VAUYTQzEfJV8Mztnl3crv2FzwQRrAiHnBTSdVBxycTIyMFaSoJwIOoE3TF5GFNiRBmLGu
lXrLchYsyn6psTMm/8s/thnWkkMlrEzCoxuRI5GUjTCzEADFQ6G7VptamVRcE/sFpGHYE5s74Q61
7zqSAxZuPqnr2NJys++4NiuGeOGgHpi2oNme086N9rmP4s4Gmfq+MWzbkG0y3xLOl3z1HY4k3X0W
WLMaDbS1WeH2yBYU42rtuoBmBgkwRSY+NhStbmLqX9SBHWFYEttzXZAz2TJDCCY+uI8wu1yizjga
HHqKMELs7ZDFJORNhQ/3aE7gQM5zhssyplOx4vsk7zEP5P/1E/A+RyVuK9P9Ebpx/ECAyM7VrkHO
pLmqew2H7w4H6aQqjMr3bLsJMnhuu8tQvxKb0ggkPP0u9EB2SV8M5hcPaRYatSHF1hd49Lgb2zJo
9O/uTXxxIfekY4NcPlUjdnI1t9zxvjw0c2f/VrBFlkMHZHw8rCbAL6yhJofge4Te8SOlcshktsVC
J3IOy7OiJ9pVXQ6qTJtfrFYnAarnuIuc9888kG5be/rnKcWUw7vMYx/KFf2Mz4eJzGoiXbZUWDNJ
8ejy1heFL3WKc2le95KB55p28pmwjEuM8lfoKjfFKIlX8mRkzUf12nIW3H4areh4KCOCt9KDksE9
UweMZCiPXHzcWhCPvOxygPIsJCo4TJIdnCbLCZqpdtyJf0kPt4qGcGDhKfP3Qapjl8g9Balex2zP
WiAQ7Q+BVr83Exd/ts2vfpnUa4rhBB2McvbgiTfC8LQ96HwsU6xfDmWokFh1FMqmy2ycObfHNgZa
Ab8JLYqRsh1uCpIRh1ssfVTtHO1HqCCjNrZ718fVAW5taR+TmUL5nTm8XypcZXTPNaXg7yzltL0v
wnK1IEtXZ8nyXNJ860y4nX69FlBI4ieGVCAY2ymC8+oXz+PsvRe2X/1x32acNSJqVjBMl3CL6gQO
nCJPWTI34sU4OQyWD+npD804LafsGDAVfNNkkjyVFsPg+TAjqS+Nxu4If8StUGnzDkA8ksAveQHI
LA1hhJk4Eez/zrqdq++Cr3ysG+25eOjVYB3ofyVNti5WYNV1y+koiYTZAWwbrMbu1V7CSPTorLo3
lrvqy35NT72q3NM1mdN0+RlzCid6NrQWhZcemE/BFf7Pv/mLM534LLaH8Fbk3czsFSKo6CbmuubT
hLHaQ/dCoRDcBw5GAyeM0Z435OYT5QjwORRZ0RBdNUD9qwxY25Stx81CisotGHK8qqMC6zj+Z6JM
AG+1ioKUcsgWp1hWHWrVBL8BAzhiNjjC2z++oZBLS4GU1i3vhrjEQOWrBWSVI3/RhMOCJqhIbNb1
Hu85akxrdrKUHqiQ4NxHrKYyU8KQ3Ecaf6i4T3JNbP7PE2WfeBjeYHbXlwEukNvEF9OKGgQyh1ST
qPyqtTZ+moTfEsLetEfnrUi6WadGim53I/qang+MAiCb8nbqUHknxYeOk/736HTYBRf+CNaXtI3l
hLogQZEZj3QYO7ditS8eO1/lPRX4KwxhIVEKh6UHlTU3knCB3LHMtxL/fa9W6FNZyA7h781ZkpCL
EQS6MaYd0Svvy57kvgWDn5fWwMw7NU4Uha0bXq5pTjVtIcHyAn3Gd3yr18IjCnmd06RZOoclB+/c
VIf7WHOkF2rxhaEiVVV9gB8lJFroTCFhWKqWcG+Td02HD3yn3DBg97uBmX5EA5qGwZt1PBbfNTfh
2rds1XuEx9u2hklWjRprz/NjXUeDlwl1W3HeihIngNdcLFbfAMqL9VkXR6FVZpdMt7JkygwjsykX
2MK5t7K8lnkvHnBs2c/dysgaJQXd5Fvr/sX6s25+qTOb697JJrVKDh7huLagGuLriB6APSb8T/VR
LkjspOA2rZE0Y4r/fmgyf7sKtmkAwTjEypiyFi7L9/xVHxJ7MC8TRJQR4mnjz6JfuZ3NRco6dsx8
AefyM3o47jKGZyNmjRV76TrgRGhDOnxB9lYXOsXARv/iSO78Bbt+lJ3KdbGPf01pKM8VxvwUabrQ
gA00ulOOSRokmGN0zdVJvOBlpp1JZ9uImJxPPT3LmWXRRjKrjuv0Wl8CfNQTqJ7U5BlOo+ebC+7t
S8pmfzg3A96Hdf5ottXrCSV1ZdTk68/E3HHsY9eeCOrUuDihoKZ5h4a1ZnPM5UnoWxxaOIK6QU7X
VXZOmniUM96FslEgKGOmIhCPqRFymkU+Xcxafo6hLtMzIQRpf/+COPvUUJKyna3aioyGIXdYQrss
UlGKYwzdH6AW1Z5oROcLlB7QdcDhb6LpvyvIL1CZTV66/d9PLy37NmHkM5mEkB6Ls8xf5pSF9qJq
mrA8r149SRIQa4JpfucuPnY+zZjaTqIURlgAmRYBFZqIr/yXmaW+zytzkTAEtqwBzrogyPQdFe9P
i8dPOtXywLo3cv05ZT4h5ao68RdLLyjTyaX/lFLPbKOP1K0V3KYOmkoqnMMDzm3qE7APmSsF5ONH
mzaD/2zKMvN0DULQHhNnfa1LtlzoVmqA/b9RBZbSgkOgNksS8g4fnmGcUlr2kVv0WRIwhtSZKw2y
bIguyV/KEfsSVfJUfLlCevkQ/IHTLIImdfnUK+8lJfNhjUq1ZCMFwOlTqqNzBk4bwPicjofpyyKd
DBpUKCnvnHf9hYXsMfgcVChlc0UhTUUiaWdOwSXAOJ/wk3LiZ2DBXFLOzWpBpTXwMkDnq8ZkE+wD
kiq2BkAqFZeXfFavHsL+utCRn0wUXmpnLWwt1aP6quYfaXXWugm9n8gYZ/KtnfQiulHqOz+8ZdSb
vU7nWUTt3Z2YYiRxPYS54/2+ALBWQsN+TKz4XDit6xtQn2g3u0pmhXyWGwzNVlnmdMjoWOjFgFFf
JzvNl22QqKfoGxo2SQbvKSqHFok3ur08LUOrd3eZeRDQFpysD3nxb9PmYHgsz8b/WqFSSwN28iao
hK8TNVH+1EfTKOvmFFRtzvc+3EeV8Nsx8B9JsBQ3lOrxGmtWknIRSJ2xUAfM7Zonuu58u8fLaVRe
0Tng0TrYbqrgT2UF5mtRB6FDOmVisYkSz0u0m/deQiHNcHMumAl154luUnBTyVTgZYHvmVE6YfaF
T1P0YPYC8OIoESPRPvYl0Hm36r39wW4vzOlGOYtlyEcSZA2iRUm0/HIlSBsktxJrVHxiM9f1nMcQ
6KGDV55KcEJvKWL2h07gQ+ZTS9djoUMqXOAhFJyhAU9dq1WJDqij4cPZfkCftfcpHXXCJUwS4C9q
Vy2kxWi0NMi9bJ+KylKHNUcffbLjXJPrY32WukqgDjRwY3FoR/8j4KqhuZQgRB66h0cg4y6evSQK
HFN5aPASgu5qWT5P1Tl9XNX1lhaprgYQOMWdNIPKMXkoJ6QqI5aRFqaAJwT88TBM/Q+NuXahGapd
HSb58jBnmzqqj/SaiYU4riCcHIp9HZbZtBGTDCGFLVJreE3jvj4L2gBptGOUcNPk7nLKfjuZh3BC
Icz4B6He7houuIG3B6WnVpuvJ9UYRUmnuZ9U1nphNRelryOqAhq3PwsC8lxoqaJytV/W3QX8b9D2
zG50uog7DcJV/QsYgFxHRBs1x9zto+cfwXeTpw84e3vLKAkwbOUJZbI1SgZ7r9uYbt9myNOE/tua
C6FgxgiFSxnz/bIMh9Nc727ieCz7EOwB8jv6PT7Waqbzvxw5CQmbp1vzazBdvey5AGVQd1Wgafp4
ueQ/AbUBnpnxxjKBqsqULnV94WDZc/N746m/zeELWh5nBstQbeJXdgjc6C8gOY7y6EznyXJJ6dgg
zsdFTmax9Bv68TnHfvCDJdTeyCTHx7lhJjOZW4fU3FAacdRQpOu45XA/SloCazLbBffgiTwIQ0n0
ZYJXbfTnBg7NCaSigiDtIDA1VI8s8xc92K51LEsxlXqGJhMv563q/N3PWZI4HHrIZkbWDFeK5s5t
RhffVscq8aTN+/FzI9MmUFzTIWVBP6sNJ+Uxfv0+Unot0KDB+gDprtBwofWIycO1y2bQZOhcHSB7
QI2QljXG71QJ2JXqqn/lTn6g+WdKwi3NmEhbCY+aNFVAJ26tTynmkE1FBROk9/HSr//PrpKDpWpu
crLfULFHCn+gvYgaxyg0N20/2jxtIel4L6ZApfPaRBzzpSH/4CxJyzVkf8vI4c9Cnm0BtixOk3Ag
DAZ/d5yjB1rXigJ93RGPsHMjUC6Vz5wXYEg6JKcCDangaCGVsSxyXRFGFWB29GNHqQr1f2gvCI4z
CCF7tzXIIlVCH4LxtIYada6aPvdGRgH4AVXBklrCrmZqwx+XbDYZDpXZcnjZ87biKIYKWFSocyCP
Ejizz/3ZafFb0jl33ABOYOArbbcrqIIhVpqb5KE3BQCBTXJwR/khlasIpVmZK8pP2zTIDkhjrdBt
R+nbXP4Sy8huuysTdBaJBtbG2TNxsRg5baYhBYHXVE3hHwTKK4yTe/rjnXxOtWoZrRtMz9oG/Tjq
a7WL7kLmLeq+xU9gBbzMwT94vssdEwrySmC01DavZMPZvMLpC8xwJZHCPxx63t+89g4+umUHwPHR
M7y0TYYPmbAI0hvpDPGCc0ZbSQv3iEN/C2I0Xc6KBHxbUerpN2rte2oiCqzMNJspyNIritcRseDO
cC1QYIEBmZoHTsvzO/TNzXA0sqwL2nr3PB4SKrbsaprQXH7wRfgTcV0hJ5rNpXw6uxVWRZatnAZG
wtjBkrENCYl9lK2YFSuGfQ+SOZzzzigY5dLPzNeQ7+WS4NiFDM0Gf0pBBfngTU3wQOvSR+E4rrrM
zg2hltYJ/tKqXmIWVeh3vrzoMUQ9oc1oWLs/qmJpmzihNzIip1FZ2UU0wnGJCt/7jP9Du9c9WQZs
WAf7Ed07jjUTkkv+rdVyuSpC5LgKyuZVDxS2COz+8SSFnGFQiXRcm47nDXbWJD7g1N/9BP4jAC6e
Kv8TvG6knasPNVpw32cgHbkI6ugx/DNjvIgBrT18xq03h7ux22tpxtEo29gBmfbmGjwS3s1DXqaD
a/DzqgOs8f4VGqyUZr5QM29PdITRzVmeVBGJRPDy/motm+6Rke++u4RICH77AHman0juV5gx+3nO
ognjLoGAtloGnOhAV4vA9vdsqTg1dfTwfrckELRsHE3MbJ9cnMS9MmcXYMnmO6WIBz0VJaAj2NE3
17kkYPFjU/Sg2iX2nK9XTuT3LCq9OhyZv1QXOH2frxqTTWV6KTPNscMFCOXvkWqNcFcItcRP8BWe
rq93YaxQdQ9G3v8QM2lgz91R9IHn0LJEbUvnFzsPKTplo5SH63JX26YRQUDQrCrexYQwgfcGdQlg
ybZU87SNK8KgnniJlUUgclTJi/FCtC03ekh2aUcFSGgCQADWCeMklopy7uAVq5n+VK0PJAiXzoY5
4vT7PWLwOkUNvPEHggEeC9qiX7eTTEqTtquvRpoxUGdbMFq9MmylnDvuxXM3+Nj4Q1NEqCSIS8Ft
3HJdBKPwDLo4HsmuV3t2KAbUzlvuEWR4ZsyBbU+htAPSEcBjoP5XCG7CrPzlIoEIUwoOb1DRLzhj
OFK6JpUMMQwTmGgX+aLg2aPpwH+t+FMVQBB96TczAmSxOn6C1uctmIc6/K22RHo6g+Hy+JYq+Skb
bWHBE9MMW+jHSBmBlnXOSk7PpYRxFoxKPSKaUkrRtu/Tl5Dqbf5ddLNqTWmuwgS3Yd1pDSXZzYJe
U05xFi0tZssTyLvn3goZrDHdKT10COtEPwDGZ2aTGIa+0XGmQXW4pSNGxjzerndPr3sdt/AqCFVh
+1ME7QK7fWElTmxx94d1xZaOu1XAy4j9wFeXYGi7cNoadWB+UBamC7lOb+Rg80MM19p19sHOW6iy
u4+JVygiZmZVgEtMHj2gOUWOn+pqh83gcWX0fuwVlru/JcaEz2/yMmvSmetCQO33cRmOZNgbRmRA
SWhuGDjhX1gb8zkUdWN3aNgxY1VrbDzJCtc1tMb2avd4h6e+alk61Qgr8rs3NQYe346ExlP3HGzz
tQlOqRNXZAs1DIXB2dozGVDWDKfWAQ67g6RYIrgXY2dK3GB46PAMlUeD73Q8BYGe2SMNKxjfq7rU
dqNZEBxJHP07EvFXIDZIy9uk73YWMQN6BQ5FTyihF2C8tqiiByDd1WHqB1uvp+N3DBPHWLHMenKQ
V+ki2aLpBPyFTOssEG+2hdBSppFw7itilV3W5VizsQVr9NdBItv9RMNS7KEr2d8LkjeufeTBhrpd
/zspfFeHQLV8qgz2aQaiTtLZWn7mh3428Rmpfi75wMAvROlX1XAhvMGabTAI6X64NElEVG7WTX1S
/wv1Xwv6SGH//00rX70UVI6yawQ19jSvJOFNRvj8sP2ML47HU8j1J2aw4jxjXDokooWAccM356Pn
wzgJ0hK5XFG09r1j8nlzssoiXlYETy48bRG+3sQe8sui4O5jrl+2dNjMh73tXfEMR7r8lGQDQFFh
8f9331XZ7cczfWfv/F2yTteYGIIkpK6hI0oYDWHTyQBs3QDWMvfhS3k4GEuikBd2YLmCcDpu+ZC/
XpvlGJMbTz4VqNuz86tDlN7S90/MWA1ZVmxFS0gQg8+V8JTmwFbJfBTr/TjGzuk6TlOteEt4T9Lx
h1Y7fSiXF10EHA5sff04ntwO+a+ZosWZOMBcdxXIuBmPZ9euDqSIJ38KqePnYUyg3JrZcoLiqz4v
ojMXjizhRzqjzu+xc5s/AnPIT1KNuKvEWjnaztrfZDDkDU+Z3wn2qorodou+WfQYQqZG2XXjzHbU
gKy2dupQ+CZFiNtj9y0NuNdYVICtWVCeAgqH0dZsKSht40y1EHBmT7JKEpBhEzaFCuXDpsTWWDS+
4bmoFklmNAZhleU9eaLmuno4ojFoyC5BkEBIL5ABsL/W4enZ3GnDI7WzZbuXy42Z+/Rp9dUrVlIq
RJzY53uI0HGELCDEiPGcftHUuh7Yzz/jk9qsUOvbV8+60NT0waIXZNV/V+roaN2RR9QbSUTFVBxp
Vi5h49RBDOvD6QEcCFgXKFF8rc7UTnH2y8PnR+AgjP43FXFsRIdlgt/0FWUZs0adtO96UyKTUSwQ
SwGaA5YtAWWMrO3hK0B8McGa71vKE6xbBcAjcXiWaXJTAqPtvA8jua0dUeTtpfEkzw4jl5pHc6dR
YR9Wz8hc8qbMJ8uEW8JMG2vna5RVm1JdJ6aHCqFdp5iL/v38OdUyD+9sHMe3zdKw0JywP9XIBTVL
/KoFZ4XxrEDGObSQrz7Ocvh6o6s3YO8WtPX7foy3LFBJxWKTmUg7HpXua+p6vYIR3H3HbAHQ3dRF
QhDiuZtP70SbbKdvDlISo7fxlQfVJ9wW6ozaEL0BEfoswVBTd6kStiPiO7NoRLnEJTnOtFpyqCwD
vIR/DNbsC4Uxieo7T+G0HwDyY8vW/lJk/OnnLTYc+BIkVwUtHcE0LFvLPB2pVLjX2mEuq49Fj3vY
LGFGxSjyEn04PbNveG7W0/KtbJP3qQbVNAnoneN1/e2q82X7dNEsjeHYsejiQi/jQLbkPoAwUDm3
RtwXhBTcDn6wUYfC3ullCmMy7/PXg6gyzf1CjYIUAQgs31cEvPEDE4Vn8wmZEB/3q77UF2cYenxW
9x2xnTM3Jixn/DGsjf5hAipiOkMLbnuQw4YAW4JtXOw2dTMOemdKY8kboUcvXkePRqIuYXjZcJjG
nVBPbFBLWtzGyb7pPsN8QyXQB/CyRTRDUENsCTV5nEug4YHrUdf85DS7rrhyyb4mQZ/aBXpi207f
YHrI9g3EKxtT2WGUK6YVHiYPVXc+4f9zcZBmZ420ksXiXoT0FM0Qzjoq7HElav2mebHImhYahF6f
HKbqGGudGeRazpq/xBsETR3xMWrHKZmnnAsftUGQthCZwDFdmiiG1aDK9oTPxmtHrZRRGSBOdlUa
d9bnlEgd/TlqTiwmklW1reyT9scmBJBazSvOkGs4UK7aXiDTLUPmVNu9xpwF3LIOzclcuw7DWwrA
F44nRqbJ1xOXlArdat9HSI5JHq9bHSQTCre5V6PcI6xZlZi0RE9TBYKhVX/H46Zyb712NXnXmW16
mfjfxP8Jxl6fF0N1etSr0bmyPoRyfPRnvbhrCFEcejM3cjxQVwC0dN3D/EFJo3TiuuBM7x4zrbXJ
MJ3dXPEH/tviHV9ShryZfFAoT2KJdFIJLh8KX9aBsZwhNaU/TyT6aTJ2/bgDAAjR58dFZ8qwQ0iT
8rQrkoWRFPuqMFGaZ+V5lBQr44s16eYTYquhLkOscSXAd/biPrGYWNsvc+rm1VHFpbrxn893gAQk
LHL++bwVIAl0iPPJYg9GosImS2bhNetGDZWjQPbOmalpsv/Ab7CDT/2CGmbCw1ob2ipo+hNydBCS
w28H0R4OvmstzBhcL8zvzm5gNTlnLMBncgX9HOdHy08Vqf8FLXkr+9Pv5xpFoXVrXrvrPpLyMAgh
ulyZ3hUIyooPFWSZOP3BobaLUtYK3CHMgDOPlropntNUMtSLHzhufUlVngZqHaP6QUZPLPVSPJ2Y
aRvqsH0RDu6XRJYrfYz2/5apmbhEEUr3SCkilscOTiJj03LcSIo9z5KaET4iDXiU8BTwCfzdAl+n
Q1fVK7N2nM9bG5JVWN9t7iDI/9xXV7aGVLaITvLranF5My2qDvTpuky4y7RK6sg4pPwxtSv6i7Ye
/Bey70LZkLi12NQ9ARtf9Sd8xPJFplI3dKD1IJ/JiJUSQaPC5UUlWL4WK9sqkRBzNU+AYw4ZXF/E
C1/IJdNLsgTz80zhEnjbA+TjmT/PY4YTDgBlhDR9cHxw313VPwC1LwxH8nG4KcyJoYKbS6vePmfU
oJXB7B+WjmIGtJ3dPaQrHYoQlgv71Jal/ZSwrEHqiFw0DNLAvSY8pE747yAvy9OJAAr42kPSjNbA
GQYYqvYPZci+M/I6eBH9mBrs1Zk0u8Pk5XKITwxXhgp5hD3UUq2BNbhVqDukTI76OTJheohAFnDG
0dst39ffLM5zNkiThypzzvVgKVfk01Q0GSCTZZG7FOKjcmiZQvV6zQlXsFJVQ7q+xywr3/b/h53y
tsDAj7xfvATJXLeyAtt2dg+fFk3YxbSXN6KsxkE4O2Ey0FH68oLkm1j5NwUG2hgRwdZ7q897kzoq
baKGBwx+tN3QO5sjzi+fKSGNfPMkzltBj9p69ux72svfhJFFqwUsCjQlIKixy+sgumCmMQUDJmlW
NgHSKA2SA8HgT+1aD3VLQRTDPdQd6479dqMP8DYBTj80mXw0oNXGUhr9Z9D7ihFoZqVo00W5CQj3
JD9QFTv6ynMNcs5LQsoB+130PB1P72mYQmV/RTQccWnsAj+2El3qxQyABIL+0asb1VlBvaD+DwV9
MUSnReSj7HcTUsp6+Uu5E31b3fwdDqjjTNDSAMoNJl8+C+r/tD14nz4vXhY55HirHjMJLYYeYdxg
BLbLsA2PU2nq/Vi2KmuVZE0XaZkHsAwCYyG91kk9hYmHL+ATChwpCQ+4CaCZM3NF0cfG4LkHwJbx
u4Wts9CPjIIy/PwDIHbIUtGFPmLXolG5Lj6BZ5XosvuGZ57m0t7so89/w0jzJZpAQaUCatqfuoFX
r1NoBVAGzAUZbu+z9O2k8XyN2ozc0GRkIET7qhu9Q+fNK/wqI/SAMZe1TGL0gFtYZby3nZbyCK8L
d1ymLd6qkxKn6JZ9s+UMidEnDCn/kr6TJXx9FxQXwzslx0oEzKkkdBU5LvXo+HfNygaI2zDILoN0
Y6E5T/QPZNzTKa4q3ngsSrLVGzOYncWNbsTTyyZRMgKghbE57HGm/ubEx8Yr3kp603C8+VjsAznz
trnNJGE587hQ06oD1Ni9KW+1FM+W6roFcx9jL98HN1c0YJISihSvwO4adnHW9WSY0f/hsvkJGO8w
YOnWuzU/aMv3pIzLW26YjN3w0/+ZsLaYbysMqNrrxpkp0+9oNkMMbivVFYfgRjEK5SEOd4KIZZf4
RI6p0vxUqVCwU7BRnD6HlqApQ8AUpuyqoYHYz6axMpkVp9s2ehhKCcxUxiMlrupccrEbJamr3jz1
twNyRiBUCG7Q3Kv/R2c/jK6Hi3cG47VjLa+mVql7fZajyNyyKy4cNPdBqqDKJhvFMhwDrK4hLGZJ
Uro5m8J3NdlzwdI0/aeXxIsHGAoI2Q0gNwO/ZBjejJQvfesE96GwYaAYN3meQ/Bu7whI7Rw1Kmmm
lnvh/Wtz5p4njpbrvoRBABexXaer/aHOaxkFQCsiVsiGs6rXvxdakmlP3wt4h7NerHY8RmA+oSvb
8A28NpWw0FpgCVEvZLUcys3hXY2/clX69T0ZKFvmd2vb4O6oTyHEcMGe+VfPtrYh03uci8HF4s/6
/hhn1gC+I7zGYH4kxrrIIjDQrLzU+X2p8LPNOKHpRet+tV/t2uwsfoeyHglhw7q0fJDlXte9H52r
GdLc4Fw09x+xrMgLQlP5PWV52tMzorMlj86U2Kl4q/82WcYNWrNTmdSPIwnn2NXK3pOIJUyko4DP
+1LT7X9k4K9qOOehW9SaMVV7AioD8oUqulwUAzcqzeA/t8CudgFHXkK04PAt/qSTbtlULYVrLXSX
KfMWYnDjptlO/cjIlmaj7YHEtAvohyRvuE32VSEeD5lqx8S9DZKmzHM39C64lVI6yjse5MJoVOZx
XIBGIrfHjcQshAihqFUHfIixO+186dOl9Jnkki31gZ7TLhH4pqdZWpkW41tStOPVG5tpe2hvnjbX
M8mMRtXVE/t6C4C5+pRZdmlqCFYZZRsOv63x+Cst/bYfzebCCnogHt0+4C3jlBPjE/wkLYNL1UdD
leH04YuB1pU6DwuRy2t2sv00sTkkV7D86CjH5LQVPg6GgCCEUJw1txVhXMUc8ipBwWaYU9nBZbqH
ZmxzYC6uzxmOnyC/a76n2R2auei+oqYYdfRTVAvgEGqWGVP5O33meF5+9lYb7UEQMcSQ6mxAaC4x
fle6Mpdrp2ZziZ0f5V4iui1G9KaOwFczI/XtDoc4ZTyhZOFgf9knFpm96DoxQM2LyC1G0u3zNeQB
SjM2HmoIx4cGe0H9+cgMScOGy31BsZ0O7aWogEneVXrWOBrQqsGUXihajZpvEoM/YBLjiFbmulkq
z/UU6EMtVRdDHTf7Q+M5Mu9rFtmgk0j1hGVnn/vSxLOTRr/sG/JiIibnjVrk/MR+iRxL6TjRLd3O
hx5JpfQeyxKX5kqcUuWgJ7QbEc7s4rxm46J6zI09e2xx73lFmZ1V7EUYzNxH6Q0gbGPV1tlwuxNT
dgiZ+evbPOPEcRbAP4xWJLqT9NLufw8mPHyOv1VAMURXj0drN+w8TFXtxlvsLF+pDQNWjZOeSFVz
86Av9VFwLcIqwOLqZ8ms4nuZsp4ot6Hm67Rsf2WpvN4SHrZc2Tan6qmjyJx1rcFsMkdlJBavJAjS
k+tz6D69d3tkJVRCcfTOJ0HEpDHGxj7eGxzEYeCeYlol6qRMffktzC2qC4ZI1U5Lxh+Zi+3xeNX0
j7eUsI8O3cyskzvmBiC7YQgXze5y0qa/hUKaGTU0ZYvmLP3AJcXWNCVIL8Y1OCUSeME8RTXALWBv
aHhdvibfUGfnqqD/5QKlm5reOrRzFFCReG1qGdwMVz0Qk3oxKEfKAooFZU9szuX6PmxbiUoX77u0
E5M12EXCGGgIv4Cov+hDsoQZnDxE2nYiYVgcpSAvRGITbuNHxXQKdjwJ1Iuc2Y6+TS+IRAcWBTpz
ja5njec1h9g0AM6PVf0ossKWpnwzDdWcetUw4+Cwp6JWC/DfdHYv1J1/s7zDkln47yWGT+aK4r+u
A09GK6wvmBImoq39dDP01NWToiGxCYim4FBJEtAqO2BtB9PtjtYx+9LjjYVd+gptiSgv0atPXaW0
8IjaVgkY6K0l2trceYO6LqmesfCjMHLr+NnhJCbSjXCn7sX3o6l4Dfvfs7svxQxRx80YoGYMO717
v1KPn3YSFIAcHau86izmVs4hSqE/NfO3oIRixAlfjM4TGqpH37dDf9eZvbaRBXHYeEKtqKLY9Sdx
6DHhHw9C48M5WKwPjMTQKB2qKOIL4Q0HeTK02Cp1w4OIn5FwMXfcNyzKUs9BrHsmleigN4oylhnk
e2dZ8RAPoaxfacokqgHFjDbAZTMb/iv7EROLztPVBeg17GmWBnehnnZLcok99GkI4DSI8CqJYQX2
jb/nIK1CIhlWhgWEsTwv1YEFRZ6Ygnbq2edpnxj/KEwSsSpTgJdOSl14Y2oGdGN6RoGlwuRmgG94
3A8qz1tKexZs+kPFR+zq1n5T6Zry8GgLeYs8JrWra8/Tiux2JnhZvk5M9X+7FozD3AHCSrdNtzN9
s43jETELeBxSw6JOcoKySxQWP8WCUUgOZl5EeXQeFk914O4nY6uiEgaW/n+r/UbLuIpKSpHa5VvM
xj1c9xbhBKJwDpz0GjHP53odG3Ghvjt5fTWbuJ8ICPkX5O0C2CJmFft+cPDxmZw867LXoJOF4kdO
yCLdBsSZd8SREAhKECFvuOrMFxfcPHnSBi7TR4dJyU1zRhKyVN8nD5hE6IStSUqTBUw/T245860F
als5aIEW25g0vQqX/V7yHBolMSS0KdRUEtHI0nIIPR933I6hL3bj4fMg3N0WvOyMDFQ1JO28RJRc
wbDpnfbYXZ5A6IBh4uLpxi8Fwkm5UczI4HoLKZI3N0Hto1NuQ9l1VuiZ78/m47qbzWXHZDo0/QyW
JV3SA/khUrwWPsflG8P0wr/AkzrukBZVvdeUH+QsSZ0+OiStQo8cAgnu77QnzeQ19QmiQu+zjvi6
KwSscrQYscNobco71D8sjnqa/3B24rxzt9taq3T9M8i3l4pgOi7QtgAQ4fBTVevvIN2s+UZjqZrP
fOS5JHy9gmznS2h1bToVTIpS0wwNN2VvqtpD55P1VfX/9fro1rthxysj9orBBgHpFm6OFJCRioNu
UI8EORMOFdxgdDRbFILd5P3W9s/skS6n8zCpCsRuH9W40F/zSO7PWa4mbZcq4BHJdf6OM8FseCAd
DBln8hUdIlBhkwpW6h6dmgj2W/JD1s7wiYpVwNl7SYOK9GvjxASH+lwAEg8CWg+q3YX//iNkj4RT
IVdQuvDE1i8EHX5EqTEbqGPxl7MRiGsjGMSyz9j5o0S6co5fyRB6ep+LrCpi+kySkSKE0Q95OVFN
C8ZiLQgaQFCzMikII2UuHSNq503QTwNWify8zEU83eCYNPYI788jlnLyBM5Hvc4KMkusscuOuBX0
x4ps6JdVOrr8bKgGmqJAvq5rbtdZhNgfUAil+33tELq3X1I/BIw+2QttRy7ePFd64g1e6NSurptH
xy+dZ5S1j5UMJx38p8fcFgrjQSc+Ex1Rl58lZ9PQ17jmqxQlbXklsJV4lGtmCmkP20UtaP7kXFQn
s3KhRDwGIoDIpC/mbqFuSeTHfXDc0vOizhw9BiwKAM0x72I5OvOfKa9wN3Nu+z4kVROXq9KOtIwm
5ZVZorrYXTQQw+K1OUs/sM9syKdlksL3CKQvMHaxFNJmQivGME5MTpvxF6QUqjeWWLdD2nmuRfxc
EW3zYVOZ29B2SvBWsyCz8CaGDI4Hco7V6MXm89041xpfMFVmOFl5+kIDaDuCNwMtIEp7iNsk+b0K
CdqYit6sTpYpLFOjfFWTnyawk93fIQ+q4MRIG2OzeYTx8PWGnhtvvFFLLvr9m1VG20s9H3D2KnYd
xnBlnxKKp6yFjMpTOoAp5xywpkII3nEeh2UtH1klN7wRb2etindtkhkaiSKHxH8UlLh5x17hYqwa
AZWiDt7IXLEfTJfV9c+JPYMe478l5plQQufjkLLNaeLxRLYt2pjAORYZYT6VudmDmzaL8hn/myuW
DYxX0iYOINoxwWN+VAtfaeXcUofKOceGNSbqIWWraKZwCqQdxTsqeetKCNbQ4sgAo3sDV43XV7Gz
E+cYMGEU2Bk5btKbpiDUoV6XxQdv56cUfQbOTzb32SxD/4D4tjcGUZEMOjOtoJSLrTyr2zf5CRnQ
jev/rLVDRs8MqEQmkbKmjySDKkCYe8GKyCEANSsEFHiUfU10ccOb/cnrwXDTCZYqse+GbQqvtUlN
GC3b553mxp/tdO0GCdV58siDhxWWcEeZkXdaZUUpCQGYj7ZrgegLK45j3qiiIBouAAsYEpq7QMZK
Mv8qLJhbAfnZbu+VLtZx2k9CgNNdB2lax6EbelblsFg1OVOoLeuXRcIlaD8VrEhp6bUnvrZ8B2FD
kJpHbbs50PUgUAIo/E2dRO3djlERCKpBHtMQ8Skqv22kqvl1Vyjrovm7uxK7983Jfy4JZ/hTvyhu
4VG1NW8i4LdpqoOD+WROQ4vLti4uZwUVWsExDEO3ZqqOqXSym85X1wH97XHcTSBX4Ab/Iime8Q9t
VgIFwRgKaxUX0SsShKtbQ6/coakb9UIGHntwMtMYOy6qBAeJMeuGm6skrr5MoELR+qOuLq69ZIrv
WwP5CHEEBXkRRJtYEA96JzvqD+rX3CxR14cT8jbkM4Lmg0OmUuUof4BEushv5NePBBHh/GfAfaNi
aScurU/pUpgqITgJA0z7U5sbbJk80MItHRM5GXQugHsKvJoZPLceBAYejSeBqkIKluZmoDlk0ODC
oDEMm7KC2Ne2SC0qx+3PautMyClb902hgaOZR4Oi/5ZhpjezoPLv08LLRaSh8VhlSZj4Xo1hKWd/
YqjRaB5iux+U0stM1MQ8CYYHAFYBb84w9ZqILKFtn1bLThPujuCOFYyKE3z69KEJ7xi7ggT8NKU0
N231GR+WPKg7yBDVufBgeRDTRHmWYl+qAkowOPsO1ZPQdzz74zGWn8AU3PhqN5D00XSrREYVEZG7
jlxycxWhgmq7g6DS2kTW1ch9NgedgT3zo7wxXsuGuJ0Nc6KPki20lgjS9ZIuwPkayVJB81h7Hntu
5Sl+g401qDIi3uECwq2dD+esTg7Xm7jh6aQuNGMXIM+Ed4C0KH3U7WnvbfSL1IMoovIorq0bV63b
dnmMMqj7iUQf2VNjSpWRiBhnEZ9AITEltFt7WzIImmcT4wypS7zjNJ3ohlVkyzPxyj1XdE9FnT4S
/+2FrkctUbADDLdUQgpAFSPoaqehPgNFw1mbtA6Z0qNjzeW5uqAwqoeR8tk3b4TJ1tuXzx96aeMy
d8LGT6hMo79GukFeULD6sRiIt1JEvS1OkdyN2jMziesdWYryBDs5jhBrvq/PozeHfAr1P7iCO9JD
O5QfGUGmWMf9KuEWPaQ3ggtMPwFkiYiV07RhIZbLb4iytFjpCKzHITygQyUxduTU0FHnSdw9PoK0
H/8+VfO63bQPv0+/DixWHZECArshP0Ttu6fbfHL2MQxiBallX/KlLwOBEPHBQJq5wDngkEOEEDYS
mT/xxneKzl+6ZOSS/I6up5LcB81lh0YXaeTTWh1B7oEiBljUIuXAfUPzNmfqxkQfeLWQno+5j1er
BViNLPvrBpT2ytY28hA5f7QZtkBP7Bgn7YLHr7AfI1IF7YJk0/pC61Xrjz7AaR/DYGPyneXMn606
o5vfVi4vtLl514NZIuq03NGDMEOP5qQu7K7r9nhUb9MPCb4ilDPoLfNHSG0Frn8H4eH36/YKnh5x
msxhpfImzuDaZLvjAZ03Hz9SOSKOojoRrlzGdRnC8L97ogtS9kuDmQtAYnKLRpdF/2ZmD4Q5UIG3
FKi8II8Ctp2YpXyd9tdtYFoIRYucdifQpNLETGnXUOElmNzLIlF73lYb/l73TfCFF8OWP2OTmWct
0EhHJ/n90Q7DLm3wb3JPkc8/ZcuQI96TdoqGFBDnflmBuqLWYj8kLBCYjrEQ3qpvNhDyvwv0BZU+
xvJ/S0By7SNUmtvBvmxxkEq3GkMywieBMKQ3ayIJrA4UMZ3Y1g3bnUPW2D/By1xQN2CkykQpsigw
xaOF32xhC9ZlmzWpANoYAvteYdKJg/gAyx/EjUCgBbi3NAps+U0BwECgy67kz1qH9a9Rb1zapg++
I7PHOjbbP7k/TxTmgdxYZCAVYtasGQaexq+4IdPMo/9aHqWIwCTfBc0ilY5I3CewiEssDRY1UrJK
6atgdz8z7mS0tJXUHvAKuosCyzXq2BFqOG+kOZkupHuFBR4Y/2xoZKPV0e6Ph5vQ/3ntvb2pP32B
QqJCXUdWO3oZaVSznBtsbUaOYkylT4iUKbbwbe/bpOvCSM+NNtQQpoUiqzPvzkQpT77JXpo9/P6b
8XWB0d5Pah28QnrhTpmxN1HaqXipWYFli8RxICQWXkUJEicaaGJAuPB8KwRg5QI8uvvR64OV6AZX
mWZbNhzmXfy0WuxQJWXyXn9Cu+vlet0dUxime2tYzg8FWtsEk9qHwEA+bNGucxaUcurN/TRVTHqk
eqdQvYcmQ5joUQ4gziSGUNklo3SWbNcvLyiy155P4QC8vbOLpTE9KmTvFdgpp7JmRI6Ccpvi8iJJ
ur4bZBxQTfK8mmOQM1TIRAkcdNeiYxvVh07Gc7ww+UM1/l5IJlGzzK7woQmg815DNr8EwuH6AHdQ
jnwXXvLZLDIhJ88pGpq4W4eqGC8gehakCJ1Q5L2yRKwmp/sSw05LEMZo6bUUC4E0l+62yL2ygSaW
ZiUwEySb1UnaRGk5cwAXiRKrwxBfD10uS6f8yEgAAT+O6D0QDKjQx8kE/+RA+RowRH4nNWDCOklR
g6QS52SCoYcYts4f6se4hslKdN3U0t1ZizaufotAuf/eS9RcODxh9y6IHTiyIkQKD6N68gld+95T
MardEaC4E7I/AeZi8blWoiJvimsucV3ovTxIom6FGD0uZlluxg5W5F2dOIW/x0xgzKUtF6PTWdtR
rowKJtdDu535YEk/z3DmRkz6teNOutjvM/FGFRufmdke/lk/STCROoLZZjMWTn8l2DGaIfqyNJNS
g9FXJtYRj3glO92uk1m+LFZl+lrtKhbJMfuBBMwZzz36/8F+AJ80Lq6CQ16EuLYLaXCLVRpkTup1
WZOO3qFwKhSYXtyzzvZQYu/rft7DKlamAoMC6UZMlsB/wK6yD0OLQUG5Cw2EQK80iuWEGNIaj/Vf
lWwksuOwJfAT/ZiDMSOI736oUpX5K0bB0P5BlRovBz3yNIqKNN8IN8kpTC8J60D7wo6N89EnmQYu
/1I9LNZPyrVOUBzJgX9B1SgcG7Ztsuiq+Elg3Q+ac3a7Qqonzu9b2xW7DXGpqGDpYPfHpNQWlHs0
VSe7d49TlhzD3rH9ewdUuBMRzDE5u12ljh0qb9NTgIjz0/X5W3F7/ZxraPuRD0fZSPNZW8hmfaMS
wtn7ysYeDbkKD6grWdGpo7sdsMeBiYgB/ao0WZZgjI06UrKovYFVHiHb9erA7K+1Wwg1s9HYB/9+
20ekayVCpjjTaiIHFuLD3XmrJGx8uCFPkuPL1BsXQ+8qo19hlvapAeQ6mzGqkZgeeA29yLAhEz5o
Ek8wHCx8KHpnV7YjfQ8WVHbbDl7jBwBUzN8CPuBx2mvLNuntfzgZS5JHfxPuFfnFlf3tuMNuOXOQ
xLruTEVjmYmyc5tjWoESZL71lez3o4er7VqN7uAf3BxYu6Fm05G2mOLTNbrrWwc23G8TrNEcgCau
hyH4FNv6qXeGnwPiYv65wyskVYGY5Tqv7IDs13VBXoLRY7kh7GSf50OKqCEFkFmT47BDLAXLq9gX
+2L3QEsBvRDGAQfRL4AyEn6HSBT2MiTUrJvhJl76h7FRAXqJanFxX7Y5+mbqVsol9RDdugT6FLfv
uNQ/ASmhhO69CB99FupMJOFh4RgkhS4+nmfmlNZAfZEP4FEaolrfXBfA3KfCMbV+zWksO4l3Rnm4
M/lgQtXCN4p/lJ732VPpQOBp7zwzn9Cy2A4Vmb8LXa7Y8MEISvmS0DF7vRmIopxgss2aKV8Tl8qH
AaTUizPr4E7y9IhuDYEc601iBn5+csgrZ4UBKgeUxnr2fOObpvZf0sn0ROjSq3fKWSwpOav/Em3+
I9B3/UemUFCwpoihhPWk1cAojLEhoWsJOB2519KE8qf/n7zSmKk+PitanUDbFM2XadEYFauDhvOB
79Oxbgu621UY8Sf1A2IwsZeL6jOwwYSSqsLjDHlEYvVkQ3FULUvYYEZDfiQY9b9USM/KQBDchz+L
ktoYIn8RfNOtRJuVViujDBjkPNod4t3Ll3nzz2WHyaNLIbclh2B9GypUQ2ZIkepoM3ZQEnRlN/CF
8KJRbwNCir7MzPuN06tN11V9fyLL5dkPLoZAsNu2soRWO6iqRrG4s6yBsg1o4cnrL9Ar+t9Bmj25
3LTR5seERLh7uQ9/RqrOGPJakIdT5ot9BTS9oia2jL5AeibymC9NPNWj49enVpblDI/D7dMlGLd+
JjNybTL7IbwA+finNtf3qrPyETwiz7Ct44ZhgCO5GkPb+SkY0JWHoLmQE9+Pw+jGaBhczUJTfIv4
B6D9NJBWqg0tYvXc8f1d3jpayUNhN7eYtmGaG4XHkltgP4WYyabZsldpYGrqYUiFBQ9zpk5M5JgQ
Bqgw9JWOwvuN/BOsYiT21NwUv7/HGrIZ+1tGV2zynUtFiVCY56taf1JkSDh9cdGrL2Xo5keVyAux
OoMgbqdd2dspKTAG+4yV/mplk73Zjku3EG/3zxn8UiM7RVvLiSxq+VyyMFNIzkL8Jsp1mSNISngT
r+8iQiCxb0cbYKgcegjVjZci+lqlKAv9cc1V26c3+WY06grJnieFXLnDW4izrw/WKrC3QI2SYEiS
MXTPEOeuOE4i34hmmRnY0br7vzZDkhmTl0BzTdQyIwaIduPObolFAa5Cw63bWNTM91wcl3uoMSIC
4MemfmmaX0nfLZgS49z8WnuF71DMS04y6xOZ20zxdOAk8aIFnj9v0CaGplnNPt47zEek3kAmZ/5E
vipth462DvSaR0liVj7umBsNNlYDMvXSDYUcMZ1Lw46aqeXf5x5cvBBc9pnvV5Bx+W814OGZBUiM
eCGG6ZtC2eK3c3nvVIHz/O11zUF21oq3LmvA0QRnRFiFc23pNRXOUOalyh+bZQzHSkwTJ0iNI9ga
1gPgiXuNRyU5ZiiNjyALcigTSGh1xNRDXKu7BLTuAJitkD3aBG3zAAKvPCfBPiVfmrgqGYE0HWN7
9StYHxIzBu4h7S0RKAw6MIeb/Lw59WCF6gNd/34oat9LE8VpL5MX0KoEAIrofjM5r+nhQCb3UbrX
zezamXxGw/tHn9JSurShyBJiPoP2lv/fIrCfQJyCWpXbxjFd59AuFvYmKKR6Xo5zzxvDHiO0Yg5h
WbQA5oVAFwpsl6wn9IsR0DFNTk4WoWqo/31ET/6U8LPrpT1mzHh8/kuK9o8BabTntU86qrggoN4n
YP6WuCoCvo223X8JUIZmjnWGDtK6Bk1oqdT4d1yxxz0oUHz0dW96s8eg+SNUWG+J4VzmDuNtNv40
MRl0utAStPygAdR+Soky8X7EejyqyheAd7lO8bybkrvv613ZBzrNVMIoSWQDzFPqjTaGSPVI1H9x
wUypZYSQ7hR42gdJqTYt1T8GcAAjxm8KWQjgd/NyoBT7F+Br82kwUnW/XfavmbH6qJliIaDnyhEf
ciFcOjvtVxfxrzCfZK8u5gU6G3VRIv12/WvbgLuaBO8OdXD8Yfy4j2EL1ehEbihGdSgpH1Pcr54L
XbnIKJDitlfPHdH1PCfopbRubncNDB1FMoROyzAcMxyy0eGFzoqbZZao6i1t7kXKrnhxEf9JEmeB
gI9OS+QzNg+dZwW5t1gh2WQ0RV3/1NwkgV/r1TC3mE63X4P7ISlFlQWB9h5VwvBVAorRDc0+3rE2
zz+jKeQHkhHp5TcDH7/pvzZQnVPlXaAdoeFDfcYUR/3HLtvQUMP+ntK1F65ot5xMWDJZdN9E+p7O
f8PzVRJy5u+HQk9/xi5x084Ux3ceh5VduaqdNs3319ux9IoblgiNO7glgfMWAruHoVl+xsGAFrQK
E670+2kJUfMO4jGJCcdq7MMqoPnXFPXogwxu2lYfl2INxHvbfAnt8oX07wTwW2EvnM0iTAhBvMb0
frE+tXXbnOcpM6063YBOroJf/vRjPRaQy6W/rfFRZZQVN/597aX1+D1KhM45nS6h0xdmq6A6n/g6
O3ZjvYD1p3Yh59WAnrbU7F9J/Wmu/MSfGmiSqTgB7uj7HMn1h8hqmE4o41kcFECS1DzLasst1QaC
zADoV3mZoWjjzc8LMZQWWa5TvlEjoPWeMAi15jTDGxTjvPwlP6dhXfQSpPrGbUut6brYd5BaQ0P0
FttU+AhDY5dc+AOTxCcGx0ZSJQ/JpKHV3XJdX086DhmVUzooJT0KkF1ZpSa3n1QFMm3hfjV7eIXz
qhKwXXQom8BfM+U227mvZAgxJKMoiu//qJOxRbeHy3ZU2WoYzfrOQgLqKxPWgY/ZoUqmb0P5scvz
70KS6ZmjMbRFd4eApd4JjemGDXyCl3fFk1r8hn3hfWgQAnwV4Nf8dooNj6gvCFZi99/Sx3yVqppk
32oz2tdzrVWeqRVldyDpWhfTAi2rGyxgB+/xfTNYHLSCYDjDtPvDTsXMD87VHWcfDmtyDW20DAbV
iQDiFlnIyu3irOsO9dB8duAWOjLrwpK9zQVtqUGG0e7q1zVLzi3SxWU8x3V+bjQyR4OKayMIOF9K
QjZxofWSOvsR0lv5DtC/AKltLKB3vj1EKN8LoI842dnkM6nd/U5WHWn6+JZThbWkpFSO8ynMsLLy
uD4QveMc+0Qvm5aLFHRJSoQEo2lWHavqdBHszlTNUUayodSbA/xN6N1raoNAEpmBib97vr+gSubu
1P0JiqFG4my+6o5B+qAmVKP8Uv38+eSae0yuKZrcwEMn8ETdvOCHjm07TmaVrFfw3v7ZsW+v/DWX
+ZcIwcQ+ExuwXTknmrpT2xcnSnQDcUSEcLhlWMDeXmFvW4d+Q+r1j0/RgZ/e9WlkXlHwCuVCLKkX
r1xHSO/F1OcMFF/J+5hSpxmhoMlR+OTc1wCv6SVqJnsQd9dSLSpl1NNSaV50ltfm96/gvqud7uX8
+3q22KgXM2eTdeh1WlegQFMOwECTwH1mSdpaauRLFRJn7aUIy5nM4227yziamee9soPwcSx4P16g
ASzdpFkoW7Gieq8Z2cVivrzD3uS0M/Kn1P2v+FjV0M51DJxNQJw2QSX8GkjiNFM/NSX6axpAF9Wz
WuF3xcbjQBHNOWQUy9XtPpwz/YgeMcDppiweGNE/nPu4bBDRN5QWBgtQam1dLBWwL0ChK7VjueH5
lfqk7j83uz2I3Ks/MW5jk1J8TJnam4TAEk0VkQoisZWMPPl4XgZapAd2EbZK9y0fYLHm6fRwNK49
332ZgpGpJ6os+ykp5imlK0OAd6TPiRh4TECspdssB4ITn9yrBwl5KilP/LOWTnrHmhtDa+1gy+/S
trfddv2bQgEReKMpEhACq2vOqFs+m3cr4M6Rhm9hQXeQr7jsI7epE4cMGGpjuhDh1Q6tvFIlWQns
UMlvEtEUzXQ1sx6aST/wyjU3+TYnE5vdRIStkttOresWhXQVz0xL8BOqcFnXaeQI5OduAUqyd90y
5QW1b3I694EDD9Gmy/y5zFWfIgRZESguVbnNVUJhFMDzuPWRvrDgS/MPu16hcGREnuuLNjaYKM8y
rAdzxh55l2Wo8p5QKBOAKCyXi96RAW46SzObgk0KhohMCOVedAqPq2psfSVrj5XtUUexuwJ8eOSN
C3K/VVBFlbu+Av3JZ3ClcXgPeGvPoPlpVOZWb6QIiyqyMqjyvUZ+I6sUkj/JOIvBeSyGc5ccAc6f
mvcQrsiQeCiDcp8XIC9Db/1ChY5T1bN+alx4H7am+82e/70n73aqV0rVDagVBFZe9Uu4y1kmz0t/
zPsuy2wyXjS//dFUpjcykrKTBf0tNAAfrOcjkTqreb0KuZaNSs4RvcJTTF7rT1J19xF9owRYqt82
cqgcq+28Mqs7l/UAsFhK3OySpYljFPIIHXle/gFtSPwALlajJnqXor5I0ffPnNSufyRtd1MQ8Iel
oqCZe9au7ZGqz5s9FfJzn00yN+01J6KKc8Rq3fZiWCrpc9RAapUx99pGcybWvwx2bq42P+BU1eR0
hXxpfbhf52Vuof8QeXupshckInDlbdCPYQHknCZpbapbgxxTHSb387xgl9r25tO1SMuV90LKx8vH
msNSjl7lQLRZmQWVj0sCOfQSA+AWpgNDdhx//pcTbkMvCTn/bkWBge8HsI+rqk/m81xdkLle+fzz
PoYEb8K8aX6CJcgdjot33cGySLGVrTGrl/8JhovU+4g7YukcASFkPOhvFp8aiF7AIvGgZTzcinog
mqji51Qa0q7I7bWXrUBDzOgNKChpVoXfoTG8cJyQ1RHF8dZyfM3jRDEFQ5fjD/v5iETKXoSnf4h3
Tcks0ur5GS+Fe3TPJbsC2prWRP7JEUUT29noiwsBcRO5Zo6t09BVnWjddO4CRkKNnHHcIQGGNns4
E3mGvsTxCI+VRZWohAQ1pRu+pyK7Do0BFDOJHyzaS8vwtvjU3VEbmD3lHR9D70HGiVKQ4g6Vscl3
5dTY5ysbYiFLzgVCkCe8Q2SFyXWnly5pbIzBPsUuyM/soiziy1p+6LboV7kiddxhASHxqfOwxNAd
BqF9XTIP356n2oWAFzDZQlyqtQ1Wnc9zcgcDVlYwqK7eISu8iI64Xwzpy9EURwkD2WrxXlDsVcDR
fHrWxMQZ4BekPzWrO0GNkVNXb+r1IKbg/oJ76eYkJ2lGXD2Lk755WyhHKlcY8atNn2Q/PnB8PgQv
o4rn+m1R9X0Fv+aPipEBxvUgT3tYpUbDKb6mGdBatyz7WLihXOcdhoqL1waUJm5spMTC2j187xxn
2pcrhBl7FVLMRT3nSh9c7ACtxQ4fxXELDgR0iKJav6ZrhvvOd4mxqRDqpHUinN9T9ABNl26MJMdP
O0hI0MuMfgpCZG5oGFOXTbq9gXTieV6NpgDBqGS++nl6G8zam/uuqOCIIVQHpBTYi2yM7cFRoSJK
NVOhEhqYSw5Xa9EvEyCxe62JRMZMHmP9NtEgg0bAN891K5IH6KXVToEdbo1zY/BCJn/L/ib2+ShQ
X9UFBF939INau6V627FcllQTxy4qQjXR+I3+3m5bu60qD3YAuj0g0++uq/ZexvDHrrrr4nJDrlje
KaQwxVjVNpEO8jo9D+vzDPmyh19Bty1c9JzhgpoypDLqEq1wRZUhuXihxbo4v/zBYe9oOlUmIiBL
Eg7pZ9lsVp5etkKyc5qNPfPENa7zBrn9r+E/HEZ5jBlqrwtFaZ2oFjzIGob2pmV5WxF/cjyWbcuA
7AekqVy/vxkNkggdHEbiFuK1K2hRwAOEoHdIEpnIXPBM0pUQZEaIm/1g+Hq97eaxZgkmkH2y3VQ/
5YZv31jBp+9DGdQg9MSIFzJAhPfkzz2WjwcPhiQ5biVKpmwNlrl7W01GP/oATvUUQZV5lZm7sY5Z
mNOMe7OYsRvTKd8OCz9wK/Qx300TrZQ+TmZrSIQU2Z+xaXdB1/KJ7OtL2TMEvHkmjUig4tJAENxX
kT2S5yQFScGUTa/+XBlMx+erpqgLllrzjiaQuIp2p1VuPSVevDSD71o79tWtTHo+z1uozIsWe7+r
I1OWcGzc81ayFLJ8AZQF1rUUrDMh2K2L9HhL2DuAuyB3klSHxC9EdHwDkUj3G8v7vpGvktMTML7T
jV+RaV9u88u5TE7lQsDGErb7cHe7dGk3hQu5GCip1tDm0MG1THVRzLm4isbd2c3VoW96HrR8dxpc
aL0W5R4vvBthHcvmng5O4N8aBg5SdjA+t/8RMzrBOrIoS/bLC/zUNGkwTinVD7nX58H/GJYy1+U1
z9ZjPjOSjBVysO7DydVqlngUJLbvKWX05lNMCRGtBmv6YqfjvbzDOAMWbOCiaxTRiHLDD2R1B5Fb
g8yZf5E5JSaE+I88sTWVzSpVT/V0CdGMl90OsMhM74hdWkugVU5Bskgt0+QpkSml0f2pfqgj3mt7
EW5cIBHKI+yBt/nEqAlgBzpoxMwJ1VuZEAS12fxkxguLSTPJk7Z29bYhKbCxqi32ZBKc6rWvNQdx
tukX79yo+QMIpI+6nZrcL9q0UTZgev4t5aHMuT8LGMctMi1tPqaRwhujft/SwPrBhY8FAirhVww0
4Ezyy/3wAeeUms3viOMwt2iTsyr1W3oj50PeO2bZuk8sQcJVzmmLYaohn1GCu55dvulD+xVrdmXN
8Ezz+ukfF9mTNDa+ZZBDkqhtxIx47CsS35v0y/B1Hz5sOMnlqBjSrblARzgnm2deuk/eLEurnSsJ
QF7NZPcb+sTfSPxJj+VP+O8jqqyHVKi1l4z2lMNA2Bba+fXXgR2w5I0xKibvrCjizngC1j/mffHh
ZkHrRg5NYCMe3VzXoAP4hVT2IkOgm9tjUju+8YhDANNMPs5jaJXC9PKp7YM7r/RW1OFhk2SCxAe3
aOEfwXERzIAFDFRHYSk9xnSnyiL1uQHAOAq2pM/Ur1nkBTu03MdihoZ/m/sE+bVTM2YWRXjWGk6O
NlbEhV7uLEr0mPdB1hdJxZEtXGZ20bXEmITGoNSvAL/fRcVVu1v3slH+gGE7tQTViUsdt9RewCbz
qBVxVUgVONG1c/6Edx6NeFowNBZ8KgIDKUMC5U2hBW22a64Pb2vKpprSMfa2zzS6ds241LXuskwU
78AQfbuowUNBhhvAhnIBFCmK9DNcacKHItOQ0nRget9c+BaSQPJMeMHMxBJk9uj1UNerQnbj059i
Okr5d9eaKBJqdhENo+bG/9reJeP/YkVmzYgi2a2zT8eLZL65JkWhoPAeunqU++L3wkLf2EtaINt2
QobBcK4kDGRXUL3GwIuFHfVg1fOs9RjSti5iDeK5NcEu3qsQtVP+HJxryVqhmVO8XD6k2CdrP9s3
VxA0hLqlD/s/1p3sjBe4eoSd0NIoaPQJxPjZc+2f1Wj7UluuL23Q4IvhqsQtRjRe8mdCpfaSFm50
UTvdXprq86Y02X9Hwxe7eb3SwWy0Y0tdl+LJeicY4yYCoBfTllHfh5WhFSrbiz2F50Rh+SyBGF2C
d6me2/6y9NYn+LImu4+EYJfD1dx6HlPia29BaKJUDMnW4W3x0txdj5qr7TtrHtnyw5NdNe1HuKYX
2SpEPKF/c2m9XbqqO9eJGUdCwwia6cFNKXI3c+zAwHQ1dTFfWsJl6YL2c3ybp/fhhhNdvicGOLFY
kNzvib3OV+uXBYLCwEbRGGaTkFHDkpD0iGJpY1Oa0u8z0zJWxt7OsInrb/5afHnHS9Wvf86KZe02
TkhzO7O54xzISUw9EK6ZuzovBHr8Ri3UslPnlbvR9m92/P90l40eBlCMBzqLBs7eBHe3lpzWnopz
0gAVFePSCfI0jvKrM+NIZ460O6hdfvpG4aa0AtrBiVgsCxIYaGBDrysjEg2J2bmc1Hb9S3fFqmxb
F9iYCyzNnMatj99hc5z2m8XoBFvp4mbB8EQxgO8JSZbRFnkd3AXhWGv4blT5gX4pSBLxNSNxTLaI
oiSVHcZvaYw8UXs+Y6MaORdr+rzQVMWYB+Z+CFNAxJOQmgWt5ccNHW/juhxWiMFHmIYEFTTEwiVq
IUPBD/LtXvwQYyY7ogbDm7Ztx+5nRMYIkImZHoZMQqPG9CPntTHmi8WA0WRG1h+rsVb8tbYDBzVx
ummtq1Zk2gQWzraX1bnTxJ8UZ+GbCT3TjyEvpz3iA6ResFRlR5d8QrXbmFH18iN+blDUFC3DWSr/
6SOXGbIP09tr2wVREZSH4PiWhMyXgSpfRNXsrYZ20rtHnscrVzd7jucQrc0YWI6EIclc2GMaT5BM
iKg18pEPQqTVbEbJCmFzJpHvfVZf/mCSs49QPVrDQQFGCfeQ1M0fl3V0G4HxEpoU1fjxQ8V8Baxj
41S0mJFeT4j2xH2aUwEd+iZyJbsDRTTDeIgmUHCVBDWUVqJFwjOSVh/T4U2e8wtTvuTZu1k766RA
RZn2D9MBzzsyJy13yT+Sl14qvtxz3fUiEDZU89qrRW0SBT2QJHFeN/oHJpIe4umdHN51Ex98FHNp
0vS+GGihfurS2okUHW0hWwtqsnOjb9JolqxjcbI6F2MKzSAuc9wDh9x2uT4RblgnGSpT2iftSGjv
ClhMz1Fgh53oUCSu+XMkUZWthTIseunEg6JpkjawNSJ4DJoMKyAqTThLXAHKCCMJ98Ku1O2zbL5C
dx3CxNVXRuqjihalwU1/KAtnEhV8AEhu10g8kqGZowQASQ7QEZZYVbc1g+TMekesU5q/NvwUgbfd
MyIH2KWMYjuWawlu88q3IwYOkzAXRIXagZi/m0qU5zPCocB0Cr4FXacJxuyYPwUA13W4OS7hKZs7
9dkNhgrEQpWMnkSX2h037xbBrB1YTJMUWFBN+N4n9DU5HIkCUmFgPXWwq/WT+D1tLPn6vDFNsVao
RBNmuC+5ccOPMzlZoXj/Zop+yDDed4RXbHbGymukP/FG82ouLIi8SAv9fuQbjC/fm1eky97bZ//d
BpiUJdgbfA8JymMAIEOJ6jpbzPOLQow1jM6dNfgdjDA7skNX2g+suS3W1ZVFx4cVV8585L6Vucsm
6G88BEejA4EwrTur9cc2MLDamR3bcBWOkeBEhFi462si28JQxwEfs0iFwkPqx48pfU6SNjIAii77
gD8UCafT7mRg+a9Nc8JZcTPWDeRX8UR38hGH9xy7Nlp3Hc+PV6+TFzfJzhJ5gpsZn0O4gZlZDG63
jt6i+5Lk4buDL91KB9JDEmbHUEk89nmBZLNn8Q5busPdv+FSfl/XebBmubURMYRLU2ofM7/B9uo3
VfrYJ22keoxr1Z+H8Z92HbPwdJBHCozdMFiZeNfZuZmkM6+xr/n5Njes/4FnGvmQWI9bY5SxKH5o
zlMi0l7sJgDf7INDtnR9F/zEn6KYe007AzD7cusN9fhGJHa5BQyCKSpgdlid8Psm818ZRaZKtnHf
oSwAP1osm8KIUuNqkSho/m6g1bZF7T0i1OWOe54yGlsXA6nwQmPMyjYTVMGfD6jbd6n3OLflfaih
kihtvJ1L1WpHcr0c5ALhkOe14SJP6KlxWaC9ALx5Bpg17dRuwIHM57Qnyb6IHzLojfKRqJzOp8iz
dVkBC8UtDyJTsQIgglVAx5EIlXg29Tb8KqKJSKtA9Qzc9gVeaZHOZ1N0dfu+sIkn4jbpOeBD/1mJ
2Eyz7vRotdCLa2wAbuQ/DXdsme1AuJprhhEk51Vn8mTyS6XlCvpfONREQZySGtwt3v8qNurbDUFf
6jTLIrmBZNJvZF20LyZE9PwlHf4U/fzM8EFpAU7L3SkK78J9hD9fz6wJCSNSAwoc5w7yK3qYTpsX
ynNRVmNUhwq+a+zG9GdpD3weHSq6tOm6t5F8yQi0ICc6JEJXyszlCCWPogRmjb5y9amDIbuWJDGz
FiFhn2bV88tNwl6lr5njP8Vve/Ktb81ns/kCuA4iOcvTNbSqxVcy2q8vHTVGYCTmMBY2PuMIwyeM
FprGjefxN0AxjjtIxkN08u9bi4HedE5jhX+voHsr2OskYRhf7xiOseFgR4HGTaMHkt1v7O0+MZJq
3rosbUorfMpZfNEjd9e0JJeJPExHYEN4u332Ng2msJ7qZT7W1HA0XOd2kiCDq2OC58J2LTKULLn0
avCzKZX5vW1GoDgozsLu7nKEZi8H1G4pcmKD3nmORPmWlp9ETH0jwBbW20jUJg8OWpmJP4ya6UTx
BHNjAvuQ5s9KDlo3DJNB2Hwb0alqbbuuYMkVus28OKrCoaRwnRnKvbMElrR+Z4pKDqQ6lAJP8XXU
5J2F8FDNB8PSshRAF34iHMqy2eYF7j82WC1eHkMwN0zY41VP4lqDoO1Q3pvCAOlJxT7A/9EDsgno
522cTo6o44ITUIKbJieBBlY9fdA1rtLh0KEGw7HVcmyS2Q3+sBHh5FExllBAsVfIeKoN8HwFeavP
S5eZrZoWH6OD+Cg0BsYj+8mVbfkP5jqlRDRFXQ3FIqmLqFXCDXrLrLVUew9WnH5ItdBO7Hw1qHog
kf4CJEjLXQxB0wqr1DZqZz8RxgiyzsYZl5xCS2Rdvi9DP10p9kkgVg/eh8NQ/EbB99fz5K2l3cc8
2pi10WfRLzXEoiLz9TOnXyiyPKmsIEhneqd6kXLOSpSlyCkZSle74IWaIPgtoBpD8s8XN7k0vkAt
rYAIpkEWXWyzKKoRn7++PzsZPgml4Xj095rsZr2VFdD5+7HoXV3H8q34OQZvLvCOOqlKNKp1MUno
UFOET5wJH3iqX3OziRJYbTqQguYW0AyiHfLC+zi7fPeuYPg6sQ41+GPk8xpLvMguxIPu0dGy4OLh
FBKwnbn7f4IzUYiVaec3aUfnv1XOViehBYA0yVYkgEsXri00V+e7UGfY/zPmwQB91Z+xOL0nN6fx
us8vqxwxqwjnBQf6YMpULFlXGW4V80XM3AIEWLxALD9WTgH7Dm7Btk7rZcAfa118pqe2DSdk0ZZG
EnxgDKX+35z3VFRvzwJh7TYk+S7dqX6z6DBc/vbm1mOqdud+U7ToaW1PRhUMrvWxgE/6e68Lze4u
jNIyEMdUmfxdh/uGph4Bgus9mdYGTnSK82nPAcGNiL8BurKKlwlXN1u6T2AUVK/6IVx8lm4uiIYl
Fvhpz1RXTHjAALmDwNoOVjgazlg3fCJRaWg/EGKzBD3FHgM2sVEmtLTQw7lzARytrR3edq1He8lb
l/s7KbRzFM1YJSf6TwO/jOHJWOUriHEoavAwXqg7rp071uuhBEHfrezS4N+irBFdm43Vcylaz7R2
Ik7KY4puIvPp+pyjrV5VQIYW9OdiYSgJaodJ2UAmpwQcRajJgxTZehL8HJhDo/TeCIb197+61/Oq
+/IIXo87J76EKDtpE8o08vKgSjFXQrkzrSMHvNXKICtRjXmZ7kaTI3kWk/jwDN1RTg4QR+ng5jG1
2w85AQgVQPIwffdY9EMzOGL3z33PFJttCn5z7YWMsaBa7W0IxQwXiV4StxotqMvsCYL0y28wOV6Z
GoI9GUjCx/ZuOyQIFrhLoRokdPINht38/OEpfGPJTUdbA0l/doDGHO7M/jgAxfPD6bO8XdL6Z1fn
en2XuSpgztn5Qsu9jLqryXEqDHOfy9QD4gZOQ999vYzAdUBCtJnjXXU80aUx0P2mm/rVj66sk0iQ
6gMreoymWhxxYzZHMKzd5lDuOD9jMlZ0u0Cm0YyTDixfdpVWFQeO0a3PExA4Zdm1+2KXL5h5jYjW
eD5WVRe7U9rEHHhjCJfmvaN+OlnnNLVA8a9m993s0OLABAAMzRZG3Hawp7gwpexqudxZRWPut3NO
rDUPK723CJQGWFuauTHaS81wgujrkPZAkmKfqeQIdSml+dbgoFIEhoWqPlEdLuQO9hzRzCnkp+9A
JMBGy3RnSdXeXTWwpx+IGRJ0tjNEiSJDBZM1r7itkkfO+sSODE1gILdzMNlVlX5j7C0Xgqb2zOF+
LndJzIWiiO8HKBizyVKzu7BeiFyviFaW74ZJVERBfnVWso0lGFvTJOmGntwKzUqRcw4WlCdvjz55
fk0LEHTqYwVPbD+aSaJC0ICyY42yDKpgRx5TJlfvxvPgVIvVLMVw62nd0hsVCPXe1pGyKBDf2NVi
RFFtkMhg4GeRZwCRrgdgxRAgKZXekAnKSA9jz06324FBkW1K2DH54SzJvQvVpxrx/Tse+ZucLF3j
20nFylNJHosExpbR7mV91rUwBT3xPmLRWccPQco/vuOqo2UKu+BVZ1hqMFpYHKKSlHyypoMVZk00
A6U5t/juT1KRTFSG1DxhNvShfyF4kybPyApZ7fWxeqNXU65nYNygTspq8WJ6ELaz82Y7+JDlJex6
A9EwwlUZkNJOdMxDO4Ajn4dz0XQKPUUmieK4yn/grxGj32lEke62meudTdZIFqJYInzauucDhDKi
aHk8fTg3cLBaJxTJzr7jKTq+rzMBGg+PV6BBg2098VsEEa/i5VZd5rJUlPRgfAH8ta3cBzu9xhhE
8Gtupi0HXB8ZyNd6Cx/akltt9M6Uc5CBnF3cEip36V38gqo/ekGv62Ysuwo2K0S4PuveLEMACYib
Y9DQZjnMyTVgSJhcOlWVK5vpxm17DqqhbHoVxZq2QHEqZvR57FTpIJwDKTYyv5EpawFIS3jKmV/3
uzZqRPcjv/sEnsZIM2JQPlDthlpW7mRjda6HAlWSS+szCiUKztgpTlSgltSmCTKp9o23zme3osG4
y6248T637KU94BMUd+UAkPMKbofRrv7gsxIhNn6HgoVK4Odn/c2XGa7hAENaV//GF9jQPrhEeWka
st+yDTLW8ozGp9EPcphTUAwLmjqvfcaa34RoSdriMA2ye0LLsSJXm9eMagsRmjgJLCGG4JM3bcn0
zGWq+rRUOo/cYZYjMUGa6Wr5QcnX204+w/AEtTUbDrpbrEGuPd8V90f3RuIOKozwyB2cEGy11Q5C
S0rwwP8E8QOAIGTiQJyMyt+/8IT4ernqPZ5LCl3VmXlSrjs8dWms1+Y6jZTFuIZTrLrOegBduY2m
YiLeoXD3RExuR5ErkqH4x28AigUShFDY9vXyjn8LdaUhG0SESapBuBeNA/pL/uO9OwhdaBKrDg5n
wIHQ6oztWeFeiF6Y49vd3t+BmlmisiTxbGKQzJOhQXnDpw5BraQnxqwJ7s4+PiXy8tJhMwWRdoQm
CZLwmOKWR8P83dbEDWOhgK8BaF1LUs60+70yZH6I6B5FbJG4qkUpqUswMT7epBClPHa35Y+dT96h
0/xYcyFqs1CY12t5+c5CktqEL+DZ8jZrDtYZpPobYjb04/2pM5jqSAXQmPcd6CQUBmx/WGdQhPnX
cR2LsuuVx4FA/WZ4JX9gybJ/XFU1EyEX5fDghsqvY5xlxnFfXNPCqD2EgyxtXmcqQ8mNC4neng5N
D0bM9fkOGcxNg7xtSIXppgyu04SSU2oZdRMSMTB6naxGrfMOIiZYdUJXHSqXTXhV/S/zjv2ePEe9
vOR6lKLfqZ4boYowABIt8LuFwNqUqulf6HCquaiZzBmY0m7Sa195XnoMukxXTVzUK7jVXKyNjvly
KJt5YHjrrwSoOHHEMqMzs94o0U67I3ENWaj1SWKgmnEKlx0uoxwO3hBA8t2lvHE6Aki43n3cBHiD
8RsFppMSfufKmA5ICQfOlgUeU+wQW//1I9U5k3YIbqtVzh8B3P3jsOL7DKukzrj+4ncNZIisUsSZ
chLmL+cp6aq5BIuU/M8UAfbKrOqOrkcNXWl9QGOMVWRkSaVzdSG4yZrwvIowB7CPPVGHSMKKHzy4
YFNNh2YEY+LAVKjQnW22KnQeTaegJAYePQPl9Vv1xFpnOleV0S+7OKQ8r0ETGJnPfzjvXl1l1LnO
DND8lYuoxO6RkoqjW3AcpX9K4or6pGzKAE9d6HBAa5Cz7jqJKlqU8NAazpMBtui1eGqk28tWrE/A
dX9lRCQ9bP+S8fVxh7cwQ4ijjRY6vKBMGurYcfAUubD+KyxREomXxcSTkm7R5JnTgbUSAw8jUcQt
UBbnjW5Dk72amjDUyLM9UPYNlQOfvlMr3rxxsoZgDEKJ9xleB94s7nErSdTZ1c1Gf5WPD371R1Ql
IrRFoY6eJYeI9ezbijFETBAr6MFBukHRdkaY371bsDg3GRB3M5ktmLJvE45UsHd6zYRQg0iU49iT
5sr6wtDK7a7ZDZ0tiHYMlXMRqdGDnYF/dae43FbvrrG6hFQ1tUJauAkVqK/RL/xiWZHD+z/Fs1ci
2iyCBPbqqwNqExvHqD3G8WQa28kJ8rWFtqpEI8+CrO861c3KEDauBc07j/YkKqejNNNqmGxtzdKx
0/vrUS667qkplJMffmsl2TXGvL6JUeqbpKqBO3lCvEdeKbrsocJZRxzzz3Ke7LIxIYhw8BGd5lJV
8j7zco7Elj5TH+y7EOInL++hUPd+1YSVNregvBstEd0toT3dfHFL6b/r/dwSHMwkIQacr+JnjkIV
NiBJq7iCnO4S5w8wvgsABrgM8ZR61Nd6cfYQdsRVz2JKVy9dRpIydMhY04eaOimL4V8DDEQlwyqY
WiGFG57lx8is65IYGOVlfk3iA0CaZ8aD06VDN+T0Esk2SYKbj3x+APQISWrypF6fxsrrwPiWlJxH
sU7g5+PQn2NDzRY2VeP2LBUBC/iPINGbjVAy59oSPS2VlfYzHZSjg34bsnpTo5v8AQn0XYodNO4G
VD80XjQyvdCNDLaGMuF3Qs7mW+bHD3W4WAAmAL7kmPV6O14l/FJxRLA+DU+/RSPS9Bxxm8gNUcBN
U7wUUuecmOupRrY8SJwSddA6khJ0N3Tmsod172cXdp4s95H8QcX/UCdgf69v5M6kwFw2ro8m4gfX
YebMjNxsQMjYrRyeLHCI+JMs1a7P+OKaOtZzX0XHbqYDNXxlVJdOhpVMA4aEadSIEf+q26k1eOak
WH9BXo5AIM18An1WVzGz5GV2pTEwjIFZbVg7uucE+AH0oh+LTaftagtdlJytVm0MfFU1yzrTDfGB
Q7tUJInDAi+npx1PA9glZTspq37Qe0bcncfQNV68FmcsH9wURYsmjwBX4q4YZfXVcaVsr9oImqrs
scUs1MbgN/5O/yn+4B1FtK6QDSsHaWT9KOO34FxegmfDKJbwEILOuY0DHDBLXTz2O+Ax74m8oE2H
LX6uVMmG7MeY4W5UWV6QAvlGjgnk1GHbVNrUW/DMR30PoU2jHZhNwgdUjSUGUiDuiL/5q7rJfgUU
zV+IvrtUpRw+Ec+h3tuXZUT55DtpfibmwsJImqhg6lSCO1LOcQF9LyRobHxhJ8FfQKKL1iCsNFaJ
fFPUkNVI5+pJPUWsxdzrJvuKPHOEHUQE2oV1l3iJNN51tzdTFj1/s7sSeJwLtmX4BsBKLaW6gnUi
IhmBFbkYkO/xIHkTJjWTmEu5olzOADuJDtqSsakYOmRXn0GziVXgysVLMbs47/ig+TVrNOj0i8U5
NrXC8tYKq5iz2asK34SMgl9cLfjE0z8EBJ5RnLZ2Nj6TQMvSWwf+NiMEFWc7fTErru2O7axWf0P2
8/9U4sAvJkD6L1zUJScouhNam3SG132dWBdPynC+/Wm5AnJY/u4cGaGYMG+7NowCh2XnrAzNdpaF
bxGMIuAFKdZ0aMMSnVxsZD84ixYHmy1b66HBrhDr6cG+3Insgl1yR3f8fqgORH+rk02lhhsE5bpK
QxVxvPxW+/f0YjQjVSA4e8BY5x/ule2i4mAvWRT+eVIULsJaIHHag+gDtge+1G5UHVX9sza/0YEp
kBHk0n+oNXkq2+ZAQ0aSLnczaf8+8eOaOGz+Cr+DKZVyvndUmanrLJEIgMywvWoeXU8o5G/tVBW5
g37yURDqvOXyf6TN/GntEeMSeyQ/Huy9OxZzdoovAqYUfkOf6dqfwSX780GOkHjkkdbr9/1rGoiI
kO6eeZTGTKtE+lGc1o55fMEEZ7nti6O6ku+xLhZcPSHBUA9dCIRfywP00fwW9Qc/9KOoHOL6vIHc
PHK860//Y3wppQtOXAU0qscnCkSyFzaRfa4sDaXZ15o5sAw2G8Uw0aHnpu4t53xB76YWb2+KbtvT
g5efx7Zz6JQPULTBzltzDQSebdzxBsYS5kggYWlwug8UmaLJ/j0gy4A9ida9/0PzQpT0WtJ8P2EK
2BnfeSHeucZZNlbRPu7Z06Q5RaBgSZ7FTzW4NMbSyCTEIIWaOdZPWBlP5u2sakK2KBv0MTTSiuaO
rGLVzHfBcyQxK4NlTHG1ddK3uuQhnPmJR0r/Nk3aE9Ae8a9zWxAJcnXOTz+ATwvQuqUL2Kk4xDfi
K2FP13LYC3hHqPRudFgLdPkaQIiMdz+R+aWEiMheA1XTNiQ6NITvVpvmfNs6PCSlFZxhs3wEgQZc
0mM1BkTe3SvKfWoc6A/1oblCxSldUYEKqjABqtI12Hf/s0+nZOmJeKNA+Dp2eAmggzLpd1rHRErr
tRZynhS+t0QC1AGRcf1QL4B3Z7hEltHzX5S9cMr7NCggvQfvQXeZbzY0gjt575kWAEA3FjNGsmtM
DuelE0sTCqPApjCGLCXvKQxB7br09k1v2Sa03csgjEEmlf9L4iQ4oFxK4AjxFORf38nd0RItuiUN
xa0Pvp2ddgbAahCKkZWHMpfvajhryqGEuomJSkS+Lo837289VerLflbzppyFaEckLL+7UsCQWJRn
QCnyJouKv2Ya0EjLSCgOC6TLD8KxiIenRev8ZqvmktETMAwVR9m14X4rTcT2e/Vb7V4wg4kChT6y
xWrR9D87emIFBjMHQ/xPA02w/NskGX2/7Yvr4eIDD4BiGRp4d17ZQQnFsy1MBh1ul9e/mJ0LY3S/
XI/ulszBF7hyilocf0YNwgZ9/wor6yPGcwfaqtMM65lJXJoXXW/2dksP92uNeUs1OmjjSrybMwoS
4nnEN7XZOPyqMJsEfEuLKXyKksHKYUt1+47Jgsb6015d0N/RnaqAexH9GaKAok0PXbn2SSt3ANGU
ALpJP1jgajAIyTSrXNJj/53QBdKoo1L4vMQyJa4ta4HG68+CkGOL2Ycs16Vvt41mXaPCambgm2P2
UBEPBUoEZm6PUIc28aje3onkSnmy9ldolLbtrI7l/YQyQnVugAU3hnk6hGiTtW9kzZ7vU7dcGvfG
1I8RxjjHcYhCgGFWeRKQW0pz/7GNpnUrhyQ1F6bfmU4xw8CGbblSVjkWtC0Xfz9QYUY4/teXF6YP
db5IkyBfYuBXmwSegykZIzFkFB6FjGywEBjxs8t/+w6BIjqscq22gqpOZYZC9A7ExgCBFRmkn6ma
ZrWxB3iL1wIkQ6Q0Mfaq7gKJZuCRBu6cxoRHRvjiDD0hOP/QnuBQqYvK5LVKDzBBxBp5CJpCH5tF
zGB2udUwo+mDBeRh3IN6p8IcaBSod7nBRFZ70ebbzbfKHEW1wqTMoruDtoR9yaJSwBT32bw6U4YN
Ho0d89C1tPGcy1CUbA9aYeJbKc1tAc+5e+x1dv5PeWsqx7/y+VCJpr2pv0z1cXn5MAmjHaYr764j
PpTrOxQY1OQSZA+n3DB4DavweyFOEmUGDqS0ToYuElOSnT2LjD5cMOqaJt8GNLkGutzpwdIIYXvj
xCcDPJv2FVjy8K34AkgIRFb7rzReEuYTy8q+apfqk0QyRO0WJlhKq7dEgT2bmPegrJrFKPSrO3wV
8Z0yWFvxKrUBFbhy8XonCN81K5VeWotLvDlngg1LSD96jmCGTF7VGnr2kb8Jvu4R2paKrAEjmwpm
B/nWbaKYP30tblLz6ah4Gjvn8r1XeH64KT4MMyA2zIbi9vgTuCsP27v2ZTbnyc5frD48q86ksJTE
UqaBhjPBV98i9d7C3pIoSMK7pdO+Ec+YScMMrMWtiI7xlmFD+KaIzHVkRXGl4hnJuiFoHy0guKpp
N30mW4tJTildgztGllC2Xrpd5+LaQnY2b1oUFwz1H4X1Cf9iv7w30NMxUd3gqIVMf2C8JnMs7WTQ
350c79OmTgQeO1t/luO2UqfdpyU/V/m5oEcJW3gPZqeUsN7KbJONWe4wMzB8DGp6dj06XRlekM4s
GTraYGvTSErRE+yA4v/qjUVbu57AkrlIKzqrVSBw8mBOrbDbGDmwMYo9TZegxRuvdhPzn2TWAXte
ZO6yCTo88oaB4rXp2saWIJ746pi6xtaVFidl01WylJUk5FlXNChxcY55xb5r0DxsPLmw+zjx6jTQ
xw+yLbpO5+mxdA2gTI73qyzmo07vGmYYVe77cpAjbp+y3k8nCIuPZZuNQfnWwKAGLce+OfIhZXxf
uSUYXxk8/U9JlPxMM+QWmZfb1Po6BgrEg791p3eC0VwhRhCuyiVtrVpL6nkzjI/X7bP9gg7b3J0M
M+/IeLolpUgkjhTYp4D39Trx8vU00d2QQSl2xrXxoITiDADn4wBMTAqYV8VjJZhRjbqeETJLKmPo
yXJ6rmqBH9cg/Me2/qhM8zehAoqAD/iAm/9lQbzDivnGbFp+uhNVCSzXpR3K2E2XWsfCoVHMWO/S
Y8Hc+SoCvH3AxJ1S1jxm0G+tsn65n9ZA67xvRBBMF7AkqQdZ6jZgs5syDmOF90nAJ8MCFujN06YQ
9wCGTuNDpB8Lufa2u1bSG6lU19lNpMoY569pNxyyCAJwo9Dy0OK9HLbRoVsBqOh6rrgwx4QxN9gv
EUuT4FRMl3BmpYWGj8VF2B48WjcR10GMKpEI5oPcs3lLdU0HJku01TpVOoNFjtZQX30Xw5R1w5Ac
fgNUXzwq0XhlK3XkGMeiR4R5PKZ4uY7PwZ4Mzh+0SxPJtQXcSsDB+SpEcRBU1uJK/fnQyLHLoaTv
FGqGPg7pZqJl4AaWO78g3kZbjnTA4NXB6r00fkg3srlHRBHfOiYTvF1Hc9vHfILGipxmKjwBzAl/
TwKlErvo1wATfSHhSfrLkuI5/Scc19rAUWZylIOlOhVFaGjP6JxsZBD4GN5gyKK4oPZy0nqIkrYe
5kHgPyeeXJFnlJr/v4W7O89n6sdbpntAR8nsBvufZXbT/6aldQUNy3XJQ2ulqbr2OwKkqW+3UYik
wGKZwzofhpLQ7PcwbsgTMqSTzoDsnXtGaeJHO8i+fl1YQS6Sl14DyiPzgiUvQqTQbYjz5cwMHYQ8
zBJ14uK2wRdgIlPFgV9FbT/tfyn62/jpg2MKpxtktYcRGCIfhpH6USeXlwriZjgyWXkfmuPlzeSJ
05k9pfyg+cTUMQUZiSomHQynhxb6xqtpQX/v9oPKz4H3IeKl1A0ucDD4dyS+hpZk2ikSqWeJoxTg
50B2w+PQs94w7IuT+xLnFdSWrdx0DR/Z83cXSYwA3LkSp4T6jh82qFUvsK3RPBWjyGWSEBpCKgMZ
+T/ZINLxNFYeHtJ2mPVCAORgvK2LvLn30fEcOVsxU2hDnGm37UTzdlgWzJlT1zapX5cHZroYhWCt
eDQJFJGsG4O58M0It7v+hem2N/1RTrKkgbM6DOWVOAvUyu2qxTJ85Wg8XgtAofLxqVN+olZLSyo1
2JPot2EPP9cr5BNhVCcPQqWs9imBzm/y/QNA+OL2dNbeTKCcDeaPpwfW/6EA2FtbbGdsLfVNrERt
1/j7eoJMXgSNx58ajRMY11wOTAGNaXiYxImMTtShBVHG7+kRE83nw074Fa+9GODkB6m5LOYkIDyN
ufxYXovAG31EQvyrW4FWlRizgwE0X49KBaN1XlYfo7j7MpQHZhEMsn1YghT9DM6TXg/3P5r+bA3r
oeJaRATVXo4xjBG3cGvqRjT0n938XTxUpQxEfdhACZFdxrdsNNR3l6LU+tpyfCq0pxqPkH4RLcv7
YbXMZnaoJzOd7+G+VC18Nal7ONFejSdoBWvnjPSAvx/KVKObEJPsOXZLpG6OUEKNzty4XoC/iOpe
EmRQuclQ0KCpPlGZxdL/uGhCDFEiwGUuJBE5w2J3WUhmQZXmvX++TQpHSGOMqxM94xxorV+hDCAs
yhjeivTFL5SRYkzRL1MiGHQZ4JaLyTxXZbEo9jXdPahiEbwUxiwMxDjcQ1zNn9TTWjEoUkfS6MMx
MR6hcRYdO5LhRxR2sWU319cSI6TkCKm4JpLrs+6mKsR8kk1xEDdYGckHQofqWa5295FxlyInOFKq
xU+EIryyMrSRlGU0IHD8SrHcnD76G+BtGQjGXkUJetOjUQ1PZgK4mrl/PM01u8OEgtLxdoudMYaY
PxKglrc/IM9bNCU20d8l4cG77saoWBNhFPHeZnGv5LjvJXKLK4eVaxu67h7rGVUGfD9FxrlQC8z0
RGGTk/9Vxlo/JMkFwR412qRPOoGgE0qxsDkX1kD6NOvwvwmc1MFNQGDvDboGuopCoXP/Q/8fMUqv
OiDr5x3tQORbO6+TctbkhD9KF/AW7E22RI4HqYyPB1n4/5DBqhongUSR+MlzscG97o7G1TPUfzrS
yvcX8nm4GfGV5MVChLpDKoWgPSx8Pw95N0jWpU56PTPbbi3Ddvd2Dy+ec7XjCf+wwjv7NwfGHriW
AJTo7Yin/i9nR39FYgfQZ6mkBxt8zuxZQdIameLhfRafXcCWxYZobIH8g9MaZH3/5xy77Mt1ZMOD
RZmocbqtgCqIGRALsHa12iLnaF4qFiGpCkAQH0bd7yehRQYoInswdQX+DeMNGR0zdJlHaXZzIIM1
DFXqU4nQbuc82vuS0XqL8y+oRY4ECwQtf/xqTsLdid7O/tCu70WtFkEC8SWJubDATcds2SXc6z/7
KIyxZnmgFk3WK41S+GdbH4h7pQHm5mJLFagHtDrwTYDeouEJZn2dNKOWhBGlli1bsvYbyaKNGqZF
zC/9avcubvOO7mjhbp7J7es38syb+BOolvR8hDo5ICwnRIRLxqlUjMb1F61bt7d4eqs+1Xmawa/f
k8N7JMMnmcGF4AXRGmwLEYx0o8WUT6SBnwO9Um6n18PsMHRXP1eHcGCpVpFJME5NPHDMFANC2bo0
BJq9P7bQhaiKjBgSaPFndV0YILSWrq25ABGKtIepOAWo7GbKbhlxbYEHA/zcl4Qu8l+TX1vgX/W8
ncLchq9vTzpC6ZHbtk7lQs37YrpVHskw2xnuCUuQDyC0nr1ORplKpArf4T1vbUNJL7L7G0wpy0ZA
6Siis/aXQ09hOor1Sb2N3EkCGO93ayFT9oPhhPT2Fc61a//kR/PW3pbmNfiGHlBMAOINfgu2f2zT
X3S1+7XriGOW+HRwgxW05ScDnTKlLaxNu+1uWt+Pe6sCnuQVURFGYANM38f8T1TvA8nqSbbNra5/
xMrTfPjEGaR93II5ww0/N8bufZLpTj3QZMBLZWTtOVuZgGSp5vNqhEu79E3jGSd+mf7b+xYfcq6h
+hEz5RgXXU3VLb6c/YYMWKLg7+pU7oxFaNAc/Nu8ovgtZ8P0RbXVsAt+PRNHPt77Mh6QvGB3FEbb
FvSUhNZ6F0XoqqrB7daXErk9gV/qos8CSsIis7FVZUKhPUAcU+Svpy3mYYa3hWoOHbg7Ch0PjAFy
zvQaoG3sESwZ6cv1grnj3xRBz1K8z/yTzegZLRmXm8ntEhxnOd8CeEF1cNc6KHT8fAi0dnVn/FpO
GLJkpnc0hjLMBZkjWX+9tf3FbKE2NrzHVMEmdbt1Bjybwq6Sc6NdYw/7+vo4WWiZKcsB+aWGDoay
SgXow/ivaqiepyc5n78WyICnIR0jz3G4iMR5gWQgCCKgFxNNwJhIo+Idg+YXimG72x1vvvPV5D1T
xzys9trEuGTAOn50VKHar9aoEjFF++XTzrefZbNFicfiNqUfPRSfWoQslCOLxP5U0aiwDLbUPlCA
hNv+ebtG/I8F06IVGoNqw/V7OPclqIiSrSwQhPGyxuSonNxqhb+5TL4jBY7KOM9T/Hz7ulvHjAIb
gfZADC8LbQKhDUWUNVrHYC262rhuy2OGLx+xUVejOEqf+eeY5P4d6N6jshaYfn0lvXVE5EJANOF2
sZntGsvC6gWDmZtlQN36dGj53xm1Zqro7P6cpD/FqMUqGyTnB6263NrOrTJX/aR1gdE7mfOSmn5X
jKeYduzVahTVBelsFz5j2UENvNzqtOOq67iLAMK6WzPn2LZmaq4aMsDexp7mNj4n+rtQvJIxizgb
TkNC9CvPOWATvPRkR+b6Mi0BgEiUEnBssqpmaqlhTMSE+eYlhS4cF5ucPxtMt0OQotHEj63U1+pA
16GI9zlZM7ugdd780BHYuohvhlFwcq/W/kqzjQfH0AHCkcRX3t3zBTQ7ViIHINDve3yF6gBytr0z
go8I6Ca2Sy4EOMooqYpXblgXoUHHtkEr26yI0DrhDOQVgAA0DZI1s1rXmGT32o27NkeqeL9g1zbZ
yDspvYFXLmQcTk8usT5SAYtgZNGzZjfYs2DJgNGSxGQumthryWpMOc1o4BhH/jRqAiQT9FylvjHQ
DWEJoMPwypybLHcvh+7fA6ZbEM10knp5IKbKQ2W61wq2wx7SInDAHokE+w2pZbsOIg40dij0LiAa
/MVk8W5l2qO7+T8VjpWW5fCuhrQfYs9o2xXs/aa99gxPvXXtMZ/XLALjlPqGbxhpC/GtZvhB/XiZ
9YmjsL2s86PIw3UMf4jreheBv4YU6mEIDghM41CAiGCiF7EpfxNWVbSGOKb6haOISU3lI9WIlHm6
q3dKEvwa1+uNn8dp7xhkB/VDXzcF7hAnd3hDqOuSijdVgEFbdr8LWHQetYPElm63fe5IH8HP+eP/
JSaVt2i/L/V1coBo8/Lq7DdaotPKOipQLgIVbSddapBGY98bF02hfqWv88b29+a5K5exOcWKpjER
zfErwfK/HBWUMKs07DHapsjf2puzPhE2mmwADuULhxQxr+i5wkpq2YKah4mXTaqVl38rO0qh0Xx/
nsOq/yBYxGzoRBpSExLkf8yl9d687Nk9xMdQ9jbt9pYg6gQIdXJUhzDfEM+1viZLsyDaE70LWgDg
QE3N5HWcFcojUFvosXncES3Kiw8Qox8UFdLqV1aK6DIqAnLY4XEgr1Rm4wbq5QPkIpM20DpSox1h
RORr8H+4L/sQVXY6mhQy4AqtCuRF7Q4C2VlVMYGpkicTZU5NUw8rMKH0zrjLY81MSDSD40PTbVcV
9WSQzie2pEMsZuD3uKbUF9ARBaUB6Z2XPuIZdCmlW7S6wUYgE7ZQyEBRLphYjn07slwHQyfopBjk
hwjfPNMEkPPs6yOxXtAbJ3eX0colixmA+ec9Alr6LS8HN65xe3SSFkks6MN28Fe98OpvDvPziXta
DgY81XPHMWS8hm94AHqJXT02nhrJNy3qvxfkECxysrnpn5H6FR7kWXvuQShMjEkzHb9OEZeUZAiy
5kOLPfdhFKpklGHjYBp9JAou7TP+MkOYjJNhIcF3lrf6cKvz9OJQua99A5OwlT20lH/kBC/VxY0I
BVkaq2sVZ5ddSBVzyuMittJP1xncr6b6tAFhYKXr+957aDnGoevUY8i49n/umkd94AFRTbNCJgIE
E0jvnkLulXNDtapT/jH9NcrtwxwvWbi4Nak9ysPwXBxi2EEUteijXanm7uG2pp5dha960AmGXsGz
LLwUSYkYoAV6QNjCUxmIGH+v3q5vNRlhuWf3Hg9RGQ0/NpZfYgOyibO8XwwTYhjTkrxCcmymvsXn
KIwICEyNbNyLqXNEVFn7gyihvY7a24g2wOgBi/WgCfU6mVa7lP00e0O7YIQvAfkUM3cnVAmKlCZz
kiJ8bnMnTdh4onNh9RsD03qw5PolHk91LuTY1rGxi2FFUF7NyxHhccTyvjC5MW7HwCd1uakrzjjw
ruGTI3NMt6rXWkg0Mc6ZG0dYi95x8uiSJjxRYVsNnRWpJj1hL0BfZJMrXFPVqYipg8pGsHCKCCIp
v8HnMgAuCFrQykgIHIXIzs/pmwagUJ3tugjjmm4w/cYMlKfy3ekzbSol9q2nyDq+XDfhjNU7FDRm
NO3dKtUmnDyrk76YXpq4Ynok/r0bI5jpwMEmGnWeaM3mLG1ykHqCphqphh2VjuIrypP4tx/hSyvD
lEM4mNsSvhPydJamkCKkcWkqEjYQ8RM6fi3XEFKJuDcenZENeR7vwgVKepbM/Q5xqPJ9YlxpfxrY
vd4MngirS8NIVKm3UsYsqKtbi65oIg4EJ7lj9MdOfWwl3AxjuvaVyK3EKxEXttHqbSHg56fMcYKe
ZHG+3UO+fBPYkdbt1MRRDGPugK7P3Y+kZioh4lLkx1TCl5mBJKwkZ6vfILFDkSF/cYMPKgiKSRr+
8BriJAP5wpN+cbrYyfpS9PK3kia4/Ia07BR1FHR/wX0Jb4WXgJONbYHSZzo2cOfletdRWehobM+G
vNHZdjSCLbkY/DtqBEkFlgaihGpyw7uK/g0C5UcSOoQgPH7d7WTC6RWBt+62hestZGJ+1oNaHt7l
89xwgWVtctJsLNBiZBKxnya6CiPvPl5jerl5KDw/DOy9yO85C87hCiE4bYhViy1WrVH6Mll6AhZg
TAadXFivzOWCRd6BgTNEoLvtmDt+15vH7nkahSXLUYnpqYMS1ZeKpPStvwipUHxgdzMw7toXpQgg
KzK+IMiYmDoo4GynUPP9wxuX7VtwExlM6GzKI/P3x4M9XPepJoZ0zZMcPKutwMKdXSXbUHlD4hZl
OdPo1yMd/vBAa+UBcqYYJ54XUGVc8smXFbYTXu70K0rvwP96k7LTuyR0NCaFmMzDoJCMNipPMUdV
SPP21I0CS42LfUhsDVk5ZgK+cvI3jmHd7jQtMnTvboEoBzBGIHbQtWyJ6dax3jWiJ3PSOqt0V+MI
p18JUokieTgvECD4vpNwkS8NbTCFPeUgXKZTNZ5NhMlqGs8KmcUFf1GsRTVfws8JWLpOXpbQ3e+I
sMpfNNW/yaflJp2bRB+U7gBqIv6fNYzobjP1cWmD+2x+M8cPFI07OrGAUkvsGy5zoqTN+LhqqkUM
hzoFILezng/q/b1oAO885qyS2+PDck8N6PBAZkvdYEt3oq6SoO1Y63dBirR/nIPKJPWj90gNDUqJ
AD7hAGq7+i15IjYP+Yv5yVEx3VDCMxKYbrre6SaLoBF5304N7TGeFwVp+M9k9VfmLB6uyVR4Y5Jf
+zICZLClmiYU0EwOlSb7bUlYLo1px/fqyxy/OrcMPdt9FOcbl9FaE5rdDtLEnIvgH9Mp8QxXcefg
tpJD2bb2DUXbUjn8OW1cC++XRym3kAoE7qp9kvIU69arE24bycDyeKLrfxeXunfnN0Vl/QJKstup
1pyCZG7f3YIzYgIGGklbxtPEziP2wIlH4sib/8fc3hKAh3r5aHgqJ0tq0f8tpNcMhDmwQwUbuttu
Zues7/NtlebcBpk2+AILBlzzyTLwjC1ghbiEdsTWaF3o+BH0T1gGDz3lj0IE7fEH7PjGKOltRfP8
98YwLuPklemtoA0IJzVHrD9zBBaZ7usOO/PPBcGrZ3rWGF5dYTed8g1aV8TjdUt1NQAYNxwLKZJ8
2gpLcdPCohrkAeIMZHc7A9ni2BhT391CBFf2l1hCo1iiRxpktwLMjaeZTk5Mrs4ukE2tw3SpHl36
rXsqN7K5yyzPi3Qwhw0ZLAH5fxZDPIeKJl/SQeQHtL0gkbkH8HrV/hZ0GB2JLRqOlhTuIT9AKXag
fsuoDAX1Bo4YSPgLVoPIJOulzxzSupaRUoqeqPLtzOd7C/5E3SQLzAi80qgxV7EkB+gPgEqBVBl7
mKLuodFYzRMT4hPpjBGygP9KvuBkgNYm423nXp+kNv04Gg6hCGbAbc6SJz1eXL9Id4+7KY335Bk1
sky/QzJ3rxc4xvsRzdEjcBVIsM2hzWJFhdjWv3FgFDh35nvGIGdVgY46IklFNQ+a2qhbKyG5baAa
Nyr4QwnNISjYl1vRWm/k6/fLhjr3hUuC9TX2146EJfKBZutmAxojRIhCEt/+yr/r0LpkIJZjT/zJ
H/FJsHJ+qUxe2TyJ9LYJWap85ANFZUuufjmLcPovbpjVDLLSv/5tDtBH4P184oAXy3ezYv5NEx0V
gFQ7PHJLusAWzyDRiShTj9/JQUEd3bjaWdxheSQgapHsi/5CSlBjSS2PKPhXCX5iDzOLH4lWD1fJ
56FOYoKRh9WMp996EfY2YCPNNpQyysnb2GH3MiPE0X5kUPOdDSOq8C0qRyDmZsKQkGm0JU60amwI
A1mTu5C8z/35mH6fipPEEn2UtDo24F1f+K21y3ltz+zaGGy+VLVYddnbOYtR9gSeI8oDxNl8ACCC
jfZyKfS60C942/s99uJnSEx+RoXI1uxWFGePligW4yWSAxBoiw1El4y03MoAE08I7oW2432wgP6Q
MpIzvhg1ilinmGMXC7YSLIaVuWYQPrJJHJG+cAV/68QNKSXy5pGr3RWB8IeUA6s4nnLBRMZ8If8V
4+zKtswScMPLNfGMpBLNeUtb5KphnikL6bc+FDBNOOluWRaBVlLlBfgVKe0LRt5VSndrbtCo40DX
5ukuvTLgVOxHYn4XVjg/ISrNP+CQiYGuqU6FopMzy8Cb3Sq7iBa6/P34KHNPE6wx0006qpmD5jZw
3707sBbpJlacLbQoHPuXnVm8uqFs5BxhPv2MaUWd9/XeMYFPlF11DpSl+p13STy1ZaY1pkFFzNEC
abAr4FfW2nhcRlOPJx6ToPp6GEh+1EJKRoyJtjYyWq0Q40He1VPzWIHAgjvJVghPavag3a9/XDNn
ZIolD07nbJ3C0zhNAGASDwCpCY8ck9eHCaxpnAusTy6N5m6fQCasQit9GedSVcR8phAry+JeEzE9
036XroNP5Rpq8AnxS7sdddhuP4WUY6aAJg665kEvjjnazqm5DUP8LeGVTx0ewLFMphwrqxWci8Xp
5dw8J4T7LOxVGt1w5oFelRe/rsSImqSVssm1cErOTgMVVJv6PMx9MNNAcyHrz020335egnB+GpBN
w7uotW9Cwt7UPP01USECzHoxFN560/bmrYbex/N+L4JTph9m6ptD3abp+JUioT9ppoA0ulXaEO2u
zzX5lKTejLK0HSPVhipd+NMm7nVfV4bjyv+1PpFh0FlsiR62QNmQGKrh4jpuHs0nimYLs8JLM6hg
Sb+DDWuvXuBzacz+RvdRGaQivgXNCgukV6vy3dsm5XA+0nmEOOSRdyRqL1QMxnY1oV8lgbfOgmKv
TQQcr2KNE6TpSfZ8gneC1MmJTZ8RPfMY5ACI1iOQ8bRKQg79CJbrL6Ga8Nwiax4fY1BpHCG/LrWt
b8irJLWKWmTaZcJ4ADfqdr7QiSX1W9j4rk8USJP5oWxZWx7qrlJtGBRhzCvCKnBzVv6ywqiVxbiO
08Y1FTEmb+I3mNSPnDkRKbXDkkgcnjx33bXUK3NlK40P1oFQe+crwCWncZGQhtS9QTx+tU3mjYSi
myNm8f3az9TKhcURvCcSr3dpmSD5XOCLEDoPXF8CnFo1bgebXioWvMV2C/4+/wDIlnP8SmwQb+XH
02ZbFByGvGX2WsoaHuP8rs4WgdRU9vWxts7lX0hLDvn8NxRAe6GCacMlEzdJqia1WNequLeke12e
QRaF3CvFs3N7eLbs3N5e6+GfN3gA4ySHDtnuJmBWEdnPIY49jKhjj/yBorvMugZ4bCCI2OTGOZq7
6Gz88L2Gli4GoQTRw39cGssMN28TeZRCBniLx3MR/oJuKdYTbr2BbpmVdkgmhq/F2rEbqqHFkFHO
OVodlh3H/x9OjBz0M1/E0XQkYgTUlCuglSVtX33hhQSbYeZnP1RwohJAlE2JDIejvUIvVqQbBDbV
0h4aCT6M9KKm4d0WttEmpEMQtB2xdHciRbMvsJvxNmnrH11TzsNV/bT9pwa5vc2u1zHH9Qszw3lI
OigYwjrJOPUESbRg2hevxeNhWMI6MgCipGQtCBBjMXDMVREI6HcTCQH3kdJ5z2NEwxVBdZcEP83A
XZzdKjTRPL9CqnNCpD7tdzP8BRORpDi0NPZLFaA9WYFGj4UY1aNOlqpp+dGsUOjtenJhGD0pBqlz
4Owsxt0vJoqAyz2RINGY3WUArxzaiQViH4I9hDy4NApsvD04t5NTz1iDLABcWkZo0FXmeNrA6N3C
C7eR8q2Jc/Y0BnMVw/w1wkVmOUT2I8XOrFU+DrDrIHKrJggTKD93FabKd3DynQHj8SP+KgJcw/Eb
tzIjh3a7JLm0/m8O/XB1+LCmN6cOe+RuUH9GOFpcIoMQfyhWtxs8m1AD2rsthMdzNuHfAMrpghD8
PMq0H77chrOsrNsVuvPn57uwCs1dIImCSU1wA/K+Pjbku9BTw+DOKLHlPLLqwXdv2lyOzcXgHjbl
Cx6aO/tse6jux1TMrsxitXpG3mLJ0AyU44IV1fVhB+X3FH1SvOubiEEEncSPY9WqVSjP8YA1cEXB
Rh0vWcQujM3o0+9Fzl88aZ5FCGQ8GQz8hSLcSWlwVhsou4JQxvR+0GkQQ3WRU3mZn9BGaXJ75jyI
UCIG75ulOnPK0UA+ohogloSQ17TJzk1iKKQ9gEI4MUqLrm6VzNzOnHmw5bLZTyXbtQZusvNydJHG
Hgh3YwRlEWfxxOuPadIBylllUlr2TKBBSVUO8yncqMSZLz6A6EgmaXpkvur2zb12rVKKmib8YqKZ
UycwjRLrp05AnN+/eRNmlcNYN/6HBaI/+qB5ALQm1qlarh9UCTkxaWHlOjX7RIXWFXjqHDXTOtCE
ovzcQtu6P15wymtXjKJhqqKlImz9tMrdvSum34J06DAglMqlKK8eOvAD9y8P+wIw/Ms95w7qktg5
6M1m1gWU1TEEp9teAOQ8gz5riSmFz5u5YMvEEsXFa9euPABjGepsHMBcYBnMRzDM2EfuiDc9KrP8
D3XSILUvP4q6ajGyYYh8hHzU2OQhjyIWu62vxMlTrsYzcH9bsWCBOIH2Rqyr1MJ2CiIIxIbXJrTl
n78UzPzrQbnsEGXS61tig266R6RuGorz/E+8paNJWdYinuMaDn5m1p2UQQBmp4w6p59lM0dg3EM1
1FEUdQCfqspU8Vc09jf1nfEz7bQ+yh6bz+JdKfd4atNUzjtiln+MEoCR1BrHAK5rg9oh/PnVQvKE
lntfz4ENZCv/oDK/L57MOA7Drw7921HvdwGS6Gq4jVgTEOYx/4Hk+ocddPaztEdCeFAsAx07Lmi9
0CsJhstOxd7EfQW74U2hxcu+LVK4yQLjhS75rR4njk14uMBnYiqft89kgJF4wqf9t6vscM850Rb+
11/MWODjrcPUoxWM4450aquELvgFHBcPS1HuwgDvRf5fbmdze+x1aP1ORHVlvT+4I7pmi+YMKx8c
cKjwrrWT39fbiH2+9a8xA9oxWjPL2krOgczSA3gHuL8Y/vF5RW/iS9Ai6dmNMMAUhRcTMdGVo5gd
yAKgz7IooYftDAuSL2nNOm8QoNAFy+qh/zs8NyuwtMExomFDeFkYAL2qbUXSgzemZBx+LK8fgby/
npn0C/tgSdpnAO7+ta0r5qd68IVe8C7T0TKF5CPzY2Dvc1aPpWtf3xy2QVb++R6TCnorxTx9n3R5
1CYDbcYaOQ0fZYedtXep4QUhJ6IMbwOKgUq6jq/pghhO/3mkv5dhMY8/T8CHqwfs63bpUZljJ0CC
Kl0JAHF06YhCEzNldGTygkW4hCIHjhuk4wAwVOhmvrBkMX+PsOqDtDQS547ZbVRXCm9P/Ut7y7te
C6m3Euy9K30sDbHXwdMFNiHZRqr8mFtES/IQgDeOKK1faNPcV7gFpdJeXUW7HD/EnZUE+jUgkD2v
yeA9gkKYyj7XX3ePbIQB9CJA7MJqpfrs93MyKhHVCVEK9NvYthNaLErx5ZvzWuKzCCPjoYpHcNuQ
nIa5CLp9zRvsXWqC2fumKyEwiS0MyVuZ/JAl+LlLNSYLtcFct2TEQrg3SfDrXhP4opmJ3rIjTZGY
FBmevsh27VO6FBLRVtXugsJ2aEdf/HXTR37HOgdZFal5rOUKKbpfVXuC0s11JiCvTUwgFNMrVJWK
7rFrntaQDQ36hAJFl9RyYBGkAXVpzJPFxGi8+p/C5g9a+g3NK4H8p8igaT4oLr37tasFQFy7p0XA
Kma8KzD4BNpA6T/aAnUsnKcIkEiOtRJGFx1td9lOyoGn6gJvO5icVXzEIqle7eGsKHHmkEfvEvX+
f/HdYTIQt05PM7bPoPKyyndHd6mDllqPsidh7652iBnaSjeCBZnT8rfRsqJNN0ffZqK6eOzYlKA0
a+2eNVX7aux5fjpU1UKEz+w/C2Is0zSqw+5voZtUNi5QQ8lIuez4q2U34ViDxMc4r9J84vBmmkQ4
voeYpYoiT8l44HvtXnnMFJEKcSHVULEGC7JCdZOGsitjoRUeL3caPCtf6NQSYHCQPOGJQ1aITl+t
Ru712yNHGTzqA94KQUNehQpPEm5NVPOeFPu88XfGgeMJAsvpH1WURfyLBRvu8xSWyxY/+O3Zfwjl
tCQ4o60oiyhsokgtRohr6+iXSkup2QCeQGrLWxU4d0hgQTWmAVHPz0LCuXer4XqOG8EmJFED1/Em
Bemkc7zWqiqUNBo9/XBWmBTnYjyEbWZyJJWyDUBAvinUklSOL9oZ8nPRdXI6+fEijD4hubTSoTLQ
FKqyKG2rJhp6xqkJQs2426v0fXYvP5RtoUuNDkzw/pC16aDo3TUHZR19LRq+GwUz+i9HUSivBWHJ
fQOX2P7QpDQ6Oj859S23Q7nlJdmfXgaZDS1ZkJBdfeug3IlkxhTpkRh5FteusRzwPkogYyObEWPp
QJJUjO1F11il2jTkTO8IHsbriAjWLMqCo3K+fLs80AE8V9+WOVIBpDoBrGiV6gl5aLPgS+Ml/6eB
9X1ug45Sl4SEgo1YHKhAzF/AbtS8t60sc99Z23OoJaL1ECnmoiciA67uAprVEV6/w9BcE4tERtsL
PbzKDUvzRteoKdxGuWKcfiRy0OT+v0BlOG65otnvkkgC48KUdL1uhGSPi9QL+BCrdZpyd147gF/d
n1wFMKczMvIqcbA/KNDoIuH6T/ggAOC8ChMgoQqwjIQYWjsnidoWCN0CgkkIrKVn2qy6o4S75FB+
sC3eJLx8rEgnNjF4vAUj2Cqv9kysMsxRRQ/4nRctHJp2hIsJ1LcLvhbF9Duzd1IakHdQ4136Mkph
lq4EZlIO8FBkW/2IwEzU8G+t02DxtMTMRNU8b7O2aSNQk3MrTlRiwomqFm3QdbKB/MFjWxM2Ea+m
Kj0lTR6pSoavuQ4tfy4ks3WvTv7DNw01ngJ4iJt2qnSYV/3i7B2iTZwttyekgqba4XhevUHTYWZ5
d30xWqL1JkAiPrq5cXgYdQtkDK7bLsSO0cvZ8mPFMb6EERmM0o0pFWucxPDYOcEtE0AX62/1gu8u
V4bNPxDUSa3L1D+WZFORMv7V6N66LyPl2usV/ZyjtOErb3zeK2sUzLAODQbi6QjIkh9CnoDluc30
K683mkBazR9ju8Stq+XjsAK5J9QeRQtv710iAzMnIa76OGk+WGLstGD4Hsmzqerwx788lhnXuY3G
vzsJF6dtyG/IvxgY183jycJWsV1qH54WFBfr8po2xr6xvEosTyGsZbvDOpyplFkIbcqMCvHB9cVz
SPmMQMgZCFQB4a9gcggib+9CBY71OCJQiKYHfrA/S0F3XQOzvY+/xgwicAMPnutXVw+XLSKPo8EA
Hmww175RunIrwKtZXbYO/H+t35mPv4ZCUkD1/H3Wz0BRuuNbvUUrXJQRoOlhnmZ0Ppq6NEZXgjsV
FkUHQ6kk2xeETK8wN9VDW3bJsNBmgI7IAYs7ChvEmaJYOLZ4uDAcBpLLhYRqeKwy6cnleo4zYXi/
SG4KC32tWhxFMvhSQSOTgZIEHjILg4FcRKXbQ5VCGD4hTExwHWDQKeRYt/D2bHK4A8clT/jio8KX
MYAub/5TvZaQXzyJeWBbNsW8y3pP6PG3qKnwk9EUj6QuB87Tc/XfPOguX/iC+EL++W6ElGffp3ax
zlljXgGsIR3vxWQbuQV8x4Fgtyp5SV4AbRlOFA0bW6yVeLtkHFshtSwrkHtKukEOMw8JB+8dkBO5
bu8BkwCf5teT97mVKu6TLTLYcOCRQhSOjVnZ29BsXRdGbNp9mbGiKNt/XVxTkcTvsdGW/rCtNkK5
f0KOAZft4n7j/6dYYcTKkm8jmmgD+vUnnf7bU9JGPV/ChO6sj3uJQMk9JEFHgw9ckXW8CY3pAQtW
1IZVoXcdP05PCReU9PbB512gPkOqYLkW9mRxq5+78ZYGz3NaO8+EgupNkM9n1u4pgl+XMSNZcKpL
UV6C5TaiA2prWxAGkwQrKrvxPUxivqnKFc0GqSvAUJtI+JRr0HIpeAaD5CSt+otFx3Uu6q+0pg2H
Q3s94UdfvisyltUPJbNaFOmHeSVnkwZZGEp6+lIIeMt05LZCAlY9Yla85uQt/fWIFIva2SrquRw4
M+Kwr2mq3Jl7/pJ8LCYgiGEeyHF6bkvPczvuy8KPRtBW3Ti+/1G2Mp6ykiKwymlPzoKYy3Iu1jzU
St2W7fc3mkRS6SAJeuOLaCikPAv/RyHAr+Ot19AftPH1LJ3yHn7yvOdz1u2hVWAsv/InRpBdjhYP
NBg+UfhSWmaqV6C1Gu1Y9aAH7V+Tm6wqS1y+iLDC+hY+v9vkHYB0YCcugO9wLDlU8UlN91VqoegW
Src8yQ7J4BJ/ZYOn/zNyFbDcYqDAq/SG83BoUwGi6C1Wezl3uRv4e9vjzysG6d7u89fQGyleNpbC
eniur16Axb9YIVF4OSAl/UiSXXDd6rrcOR+sIKgMsm7iiG3dAramxwesSrkOaiffcLDSdW1LU6XH
mTCOw4stWcD8Y0qcH//PZhk3A+0B5Q4qQ3yBefE2Mt5oNL3kHCHGH40vBWSYBZk5AHIu9fNaOg3N
+/cgtWxm3gkVsAQ6y0+ofqIYnKD/RHuI2P/4qu9dISR6CuySZEP2BibibZ81Cp7blHq7OhU5rDdg
jylwioXdwc9LyDkWcpYyV4pX663NqWyW/4UcBR9QpI9JoKS7Tacnlw963DVZnHqHqjyZhi68t1/C
6KsYOC9qGv4nclS1WwNkpErXLj4ls30BvQjhb/ZX6EYnUUakc489B1A/5vdbdTCxZghKgX08oqoM
vJ7k7y1dGhk54aCjtB+aYPCMEWUjaWwuc/DV2kt/6bvHhAm6Ll1oJa/MjxgQEd+8k8lblWgfiCb6
po7wpv/X9AzY1gFrTfbI9sZj6nmDN/ooAtowWb7COUxfBGolOaAvcrc+dV22oA4Y0awFeAayi42a
Pv8fhOvLMFSeZoj3OdiGCRLltpR7rjVCHj8OJ9zFMjvqp0+qk8EgRuekxpRM79VhS0VdD5c3yhN2
kKIZdWNAw88ELqivIltgbcJglUgFqBs91tcfBU1L0EBJKlDZrOpvXVNXcvK2rmPWlkOdXWPAMtn0
aekO4rGcm5d7NrSd2Vpaksrls1luB35Ym7GByCgI1Sl7v27r3inMWOJs7utW6aOPVN09uwkd4tum
qNgh5DguWLDDEWD7MUovYB0zTLbL65oTUCBtq/+O4FOdT5JNwbasIY4+HVofjkEjkyZCrbLOv50p
1YVz880yavgbHInpQB2hW+DSBcz6yItogS6WwasfGujkVZE5q6shSP8M2b33VYMceL3+syUSjQYz
boeXOxV9p/4MRzvLVjxj/CkipyyK7yT5M3rxEuWf3+/D0m0b3XsrZ3YrR0PUHTlbGnrQZ/9P2TH2
FgKzalIfB0IUxJC0TZCOaH8ZgkvoFycvY+ID2zvw2fxA/XsUF3G+q+XQ/VhaxBPQrbpwNxHORPtP
S7ceLuMfl7T+mdWCSJK5IEDyXYZ+lJ2Jdd8NLEZ3TQom42GOnmuAaGkFkNgvWqiPZtD9YtOnD/0N
K1NHYk0hFeeHZTPvUPBTyuIcLdB8NGunwIL2WgAbLOWNFLVEHg4A4YhSrDrJ1jmCk1MhNN9BOIvV
/gViEf5RP3xfuaLkzIt9ObNlm4Lm1zNWeLAY8+ozbnLRCiyIdO8W1op2IZZ4uksbnUh7DqxGFbO9
hF8SZ15mjKr+LJjEz1sxpNOTe6+osjz7BDQSl4LMNvzpEhDz8z8yW9t5lA4Ha81t1FVUbM/yZ9Rd
3vfiT4sCgAIAeFkfUryU8T8+VgcUb859EI66bIZZmGeCn0MMGOIZitydh2xu3mxPPdV6XYA6Xmd1
AtPSNrraf2mwgtoXC5TLQ5r6Ef9YyR8fUhgUgpka6smMF8balCRjCkimm08wYTvSvlCXbIBfJsjX
kSf6r+ROXFe2vi8vd5naUw8o/tvmJ0VzPvnBFUdOy3/X063NB13Z4urh0JZZSwJ+aUWSAnGw3AMg
IGsADt/I7ShcjYZmPhq4y/8eogcbI8pf+flNgCblL21xz0qKCKt5qIVtOdfIy3IpLNpzssGhLhl5
RurnVuBKkQnoDQQtrXaegyrUhX9ryaNp5EUAq11IFny4PpFu5P+TfwOKIvKk8ehOuhlBqfTf0GEE
5SrFpNvAlEmLK4CbnC8ws0QpZaoo+m0PnhEuJTv+VkSOtJly+tUFjZO8R0UUxZYd52HSyL8MpcDf
Z8HKkvazCj47t62uuqaSzJnGem4RBlONe7mCq+7JuFmYZDfn6q6sgFvG1j13STNKxp+AdcOFr2ij
OZDC5eMFwu0pR/G3AxuPNPpE0XEChbBDqXfp8fMkv1ssGo/EIjwwHbjMa+op/KHUfSiNdNCUrZFq
nP1jYHKvm+FruKklFTCkQ6x2me85D0bVxF5lywQcMPGkNAiPOGNIJ3ljEw5SXYE9a+4aJZlKOtsi
Ut1sQPE0wzOTpP8JoOasAY5rOZJiUiIQvnXICq1ZvD3t7miKBzhzvJ01ZjHdMek4mVdWXvLE23xW
gt7hMKo1FSDGpHnltO3W0YOPV+xkzx1t7DvtF7+OUt2PbQpjqOZqvol7aQhM7Hpi/RDz5qWAdgS8
gxpaz4WJjqyfRFEysaZPB1I958c/XBlFOaou+mgqFxkkazZkRez2hPmPtoSCzrHZs4cTjjB/+/Yv
OpRMKf2iz+CeCnIpbTtDLYWj2Img5279m+9NBcjUmfgTomhSSbmSOCkt44dICRyipNdUjlbBRin2
j9drOzBdwDEnuOCUGjQnGBtskVFDWtqUS9H5FA6cLLzh/9TyvQ/W/VNYQPzQlcT2uiCtdM23GSvO
iyOj9m98eS34qh1u/IQ8b6P7ZGnZFyG0VkyY5+myfsYvFmuvUutrYdFxtaPrbQEpaEnhGwXwo+V6
nxT4e9v7PLV87Lv8545iFv5crk2nZ8cHMbh1qcMu0HHGrcrEAswxOnGT2Gc2PsIOf126IpqYIoFc
acpf9DOVCJb5ynplM6CU0yxO7OofQ2ROWpfGT1Wv3hqZ1BXaGqwBaR9KIQpZIZVR/lQXZ/ytHcCj
vqI8ePeNSjMQgYPQ8/HIg9J11WrpoGtBcoKpzmh5W2pyJr9FkSgxkOMYbAl/MMWNoQ06p1Xy5GfM
2IRe3Dzk0gw2VaOysiUuU6FOzOd3nWYIhocJl7/ZurEn+qGxI7ZkgVw8+Knrk/NCpSD6g0dYuAJR
KN76QDsKbzOZExPZGosDmLRZ6ggXD0Qn3XZuR+60m9VZYq+CCtxD91w7nynnsYdeskNNe9hboBsp
DFgXvrXVJr3GyCQiuQ1AJCAAti22v5YX9ZbIPI8D+cG72SYAkDik5ryISLoBwUogZa4jbOP8m2Y0
o8pGOD0CR8Mby9wOJVoB1Cg+76x5p78kTk5HYndOTtBsxYOZKeZB2kgmo8AYw0IXJv7NBuUo+TN7
kLbkNmhPkF7DzOfrmlE97qn43K8DQtmlS7jL4DulgcxsBA0kmlj4aQPBimR4Id5ga0xfpEVkAIno
u0dHIEwc8gGCbXQi3S8G1QDI5f7/w0HlgAEjQ0QqaN6Mas0xa+a7SoWOJ98FOQDpBOqerb4R7lgy
3cl8llb+Pk6o0r5trp65kxmyhBRDOw34tOI42Vkypg8WXWUHiGEU4ul2vyFkiWfdFqCbO9rw8jmd
ILGsQH1f/CdFOcBVpfJP1GzOFrQA4dudVHXWmXuKw0V4FTVDy+q+/zc3WStXZZOmGVfO6BnVOUct
gPXVsT84NRWFeQWoYC5/bXVYg/KNDyhzMfPFNVvgG9gEVHZmEP+wjZ7+kpq/E0Hqh7A3VwF+lx7c
byKKi13lKNaz8ydy0TzdQB1rC7sMihMFX+td0f3oE/zGY5m7CteOH331Mjgtcj5zSZeM0HzJel4u
GaEP/BKHEvEHAddo2/hn0d09DVzvTkGomaFqJg1NkC0qcCCfawTSZz/qx4a9Epw2DjL9+A29YBlo
zz2cuaRTaU3iZ16rX20l5kdi1Pbsf0xwdzEbBTf2Ili4NyzEJ4U5Zu7IHBcLT3L8d5snBu6R+uZ1
B0gZgTHBlHwmCZreiqtz/Yg8+O3Smsyt0j/75IGgN9GGA7GdtQ+ACwwNRdHQCJCyS4qvv7sYDT1D
k7A9e7+voLjPulekLoO/eBE6szgHLS3NsmvK1U17fjzTKtlrU3fuDBcxensYcfjeN2czUh2DdAhJ
0BbdFXIDcnh3J4C5z8Jv9AkKziS5li2oqsgbuPQetGE0iAApt0kz8gLN0aGLz85szdHQWTS+QbJL
P8hBIo8HDYzKOp/iN9Tm7A+uSgOMGe9g1W3YHJMH4bM/nDYSW7PqsKQtGsiY0GLPJgUQiBtkn3An
FOS/R7H1X8NwPcgHGTsc6OJDq7a3EC25TGcySz0bTFV7SoVC0O24Et+A0I8GcC5NGf4Y9AEGnN6s
6xw7d50TKRewtrGsphcB1UqmUilU4dQ0g7Kqs6IK97spLHlF7vpzxO7wOkFXx5z9liya4GJV+nAw
s0kvoIN0GcfC6cFy2lJYzJErx0IcCuNdg12lhJOl/6TNBBSSxOcRrxVWDkCJdw2TpeKVZJUAlccU
6Z8O8C1uAna7DgU/60Nvq5fUQKhiMpfka1627OO2kzmw31ENgnc0ph/7OdqD/rga9bahE98L2n4h
qn8L97b96yYt5a/AT1fzgH3b4ehk/qoZ0KLXzwhWBAKCepzY5FQ3t6aqS+sCvmeageawbq7r+ofD
xm1uC45veAFcs2JzczE9X+Mac8vnymG759GDxgrmHsHF0hWCZR5THbjtMjamGTsus5ZjhSrdw/AU
FOguX9jePwu3JyixbGZct5LOOI/Y9uPgMLWXuclcTdkuIFiKUxNpGmx3GdbNBXzHP8mKtII+pzag
Ar5Qd54EfNaC2SMScvAOd5XOOvIzSG6kU5H3KKPdwC7DJg2MRm01P+wIdbITUOfryJF5MdCk/M1b
R2P9RUGJ+VOgSqWNZTlKOJqB2NvOaXSxGolJd5Kmqv0SuBWZbyN4Y0YJjMM/G08vDY7VKVDHhLfc
OyJcSvwKWlwGneXJz6HNoYbPa/dKsoTn/4/ji+foRL8asaOeonwlRJJovqExKB3cBYkTAkWPGWNW
84ht32AbNvflklzbbKtf6/hRQwETo1IQv4C3TesVoIqq4bh2rwhOytRCSiJTNWpzVpGExuoChM4p
cGEcMKzm3gtEfp1JcVGKOQ66l9CWoaGUvO8vAvd5eMz0AX0q8+9KpfM+P/rlcx1Z1YgDyS4WU0n2
z3CXEoA4L986VsbRGiuuiwxP9h+3rqiAoKLeUxDXj/zNF47FAdHF6tlt6csYen5x9giRC8Aev+tk
PgGYohIyD20cAOLWXW0cQzZNUn75iMHDlRFFF8B+vcS/FxfRg8lxxEeBIFw/CzSqzJwHL7rQu9cR
wYR2YR7I3wTDayz96ATctLSN62ylHypaAan5/81ifkAeW/yn7cYtRFfFDWJk8VI+teVsuk4Y4UW2
vxA/cjsTP8Um5rzDrFsOcPXrKY06TBDH3NRlgMwPOEACAugkaImc6EMduv/BFwZz5aYeZnwAl5XU
dGvxIbL9LaJXH+tgreUMg4sm7yxK4uzQzHhsesv7tZXjXYnQ4q0dcJhaKT73lCH5QDSPRc+IL5ux
J+MQQG81y/ZB6LYtjIfX8oT6GbVXiIxI9r0X7lbmB2fLeDXDf8ivO3MUQXr/diDsHgEucVUUdw9V
2IvKR28Jw/Qh+d2W1sEIDyuoECRE1kFBo7UYDpMjcqdZD1E1l1kgVF5J8qH0QyLv8wb4Q57FaaKO
rmcsGR0PzUkiIk3qJ1Z+iNcjUfPfpI94/p7SzFLrfykYo3OUTgF5mq7AsaxMP0vHMKC2Dn7yeizd
DXY4uiV1u3SumcAo+HBp19RwtDc+5UpGsDxyzMQLd2MmRJbglnFSX86f2ZcTiuoEOaiPXik7CZko
thPwMvHV5Js8BDfnYY/6McgIpuTbjIJDv7e8Rf1WM5/LOQzA6xQYHavhe3WhZVJl4fNcImNnLoL2
u1L2dXkYoIzFpb88RRsgWyK5WB3uLxVAi8Anq/Epx1eOhjsqI5hmfX+m7J+0HpebyH6z4QMeqKJF
PSSMGmwbX7taRpllzLR+ejbwWuTG2yZ3uRpeV0jPnjO3basQ26gYzgx9EPiP9OoV9T0PPWsvncqB
DhlCU3NmcxXDMR/kq5xszUD9j32XYqInhvyCPs3eS6y5a1H/LTGJCqR09BZKZKMGjgjyQ4gTGDof
0dsExQgPW6axd/pUbS+2UemgjCLC/MBw3tXPp9803DnJC2fB7N+XEqMgJtbU6GpMspFp+DdYJP1v
WRn0MvOBMg4st97i4T0MautWaqEZO3RiRsXRQLQFYEEUliN4Vt5CD2GHloQiRyeUceYXiyyW/a8k
M7RzJO3RKXFl8Y2hk4JbogDxQZqLvGHsA4Ldn8IWvspiiuTKYMYbXNg/MEEe/6D2om+86V1bmTdp
pe04OSgbmwaT51dj9qCTYEZl463J34FN02UYn4ES3rN+Xw2S3Wd+ZRDg+U8MwRW0YQHU6vaf9BvB
oC4EfZsuJ+WLdtfYIERPtiEIJb+N7k44P1cAAgG09MEqKIStBt3FYUyvcB3snPBEbs8r+4qxhQqw
B1IIgzM+kOJ6LuUP2BkoVlD2sCFfqdM9xEkW5uoE9vkGIclmMMl3yJnxjmFNAKjwbz1teoOOTqt4
Wu3sOt5PbMg9PuVunNN/XdUG4g5JHiTVFNHNLT0wAb+FnRLYW0Gf5zAWlUEkllGyc+/5HwzslHLf
LQqEzGVLgvW80Mev9nUC+2ff4UnY57MuHPa6RtfsLG44bVnyVlY8k/kRUnvtA64D2iRe11Or60tw
IUy3O8MfU02NX+kMKLrEEak14SN6o/ptWEhszDVATr867Us3kECFk8XxUFlWuoZwhN0ua3DKPXWK
A7fh7LpR0XY/XWToU71ZSKm7Gl2jkcXBHj8+gZwbKtNYZUhsWp4Q/A9XidrfR5xthZ3o98R6NncU
rakahPevSLhvPkLtdbCE/z/pSfGWCE4bbnN4JsHHvU9Nq2jUMMjTxgxbar3/iwgD45dQ99ReDzLd
+c6bz3BTq51YOFR1NfUqTyyC+lQjbkbIUo15WdvTmnMOCQl+iX8p0UP5sNckScfWQtG+E6f9Amz/
RHOPtjCg2C32bNYNVrmxes/w/p/pyZ4Tv0CLwXO7W7Vej7Ul5YP5FSXT1CAtg/rbFmoAjJ8eP8KY
pOb0JpDuupTLycBfTfceTgBjg1gDnYhlmpnUvDaVN4oWQVcSaOnEiDm2p+i5VukAalhS9K9cZLFf
gS81H1YeJZyLUIbyKYLFOzLF5IwjCisWdA+ZZjlDZiR6+y1FDPUHNlcz8frG7WiBCb8xPT5PbEMF
/dUw3SojvNMCgE3lDK1DNV/PsIF+i3WAFJe4NeqHBIMmgJ/6LJdahHlOwOJkLF0S3KAfw9DcT6L9
CRl7/x3m4t01LMR4y2uyO/Oni/kGoRYnE5yg6R9eNnyXbFJAlwNTKRslvzm70CObse8hBPSzJs5z
ZXpRmZeGA4vr3bhOVhrD1J06o0tgux19qPr5opXEKttX1emo26Zn6DKfUgeFLAaE+t6LbtXUJGtA
ICxYcePwzzJpprTtYdtLyt7D3BPgwrafztOtiKNfAVTnGBblINmt0ABx8phP25W4dtWocAMBqhcu
WuItOCFkvdsBf7/NvoG/Ll0MPCy9RU77Hbh/5Lke82zDTxKWbln5+mC392ca3eYvM0R/7PjEmP/T
2ZwjdgmUlx0Imn9NlsW7i6nrrlMtopuWapVtMSxO3galdgrJhtd5DW6xp+0ebLp9JqXylB20ZJ2k
QenSQzvBKIWI6PcjVQ5G+E/8QJ1e2vB5Q+3zIJYewf8aNb0+eYs9Ddvh2gWrozheonhnHxLfAOAW
4rIu3Ssh6VJ2f/vwxiPUVG9EsKRYNk9gWQw3Ke9eF8GjKxDNKLt6p2sPF2tbUrEONGDDuI7BcrfU
Xhukps4/UGOoBPz5n1vXZhyvtnPYALhyOkQ/eRJTaKWPeIdv+D1xDYrLbv//+CGesWA2cx2SQi2N
GOBBkH6Ft0TJuKh69gIjktDCyULTVLtoSy4flFmRFMbXzhTtMuLjwJ1euFVCF1gGcFt+CqDxSqQB
OHjJcmoLuR7JzAN+N4dTzGS52h0G+Bse39kY4Z2w9W0/mdjLydyMaGTMf33NgpuD8JGmJZ69RBB+
osqgEg29eYJZq9yqGzyQghNp7o8Dd7v4TlxJZJqccyl24pFSNmcYyvkqrPd4iu/F9UpqpSuK5fT+
QhKshKiV5NNrBtG+AhsS/lRW/7srRkpjBrA1F2fjhewm4S9mNKHysfAOuHMjppc4cXpduFZZ9VqK
efBHadBCO+0/WsJscroSlVh/Doz4GCNMxb/Arj8UjDavIZD8+xfs3/ONMywKLsHBilyPjeAYAk+Y
Y4HCBzhia1gqHrq3/JVsmujSLSMt7NSv7YnGZIFZR9FIbqcBvn+ZNuTqaJ4FxteXr+vbmwS7ovW8
Jq24Ovsa+jQ5b9u6/ClU0GTQa2nQOFF2IkApwhDg7PFMkT0Ah+BX2wpvOvKwEU7scnymdK+XMBoR
6YDidIXIwwQMjT9UPDtZHG0Kpjt7pEuwYcAcmTnzFCZDZCALjcBRRcJU1WzkbGYJeu5REwJXwTqy
IOyQDaxj8ijUY/9dhmdq/mL03Ajc5ydjsWjIDAWSBgc2u3ohLB8OPBFN212msDzSQ4Z/gcb1tYSB
OX2TyDKCC/RQGLy5izTJtz13gWnlH2gytOjrQ/r/pTQxXgStCINSwR7nNcSFlBzIhbvOySXSl3Md
ARc3gtZ5PqPNh9dBLIOp0MEbRGNhk/NPgKvtiec/UwPyF96GFBoiq5JtYEB5enaxZGgjgIWIP8+C
cArVF0z41Gyk4JoEOPLhZkCVz3XMOTWGey0ExDUqYqZEMo+XyQ7t9IHSLCIWQojGZjz+nxRYQI2R
Ya+Y+xDmeKHYox5GvXAuvBWMWpDtsqLRI+Aa40nB+4yqcCnreHhdxw/uvRSSasG7bBcmVZnp7EDG
s1II28v2KgD2JAxeCOC8TN8W5XJBE88GNGaYjnGB+wEF5iVCM1w6IvQ6u7+1q0whCbm1Tq9wQ7/7
0V8EkTMUP+y6qW+MrzDQHFcDRPKzkyE/yIPuM1HHgSU2hidfnSmbgLXuB1CvE2TGp3RaeGOIUbYo
VsCtysF852Wqiyh19IwCwxL/1059ZBDus/K2PEKkfGUCudLIpwdmKbM0cY8imrmVeHSoilthnmCZ
UsdoASg3/plFTuVoUVpCO6YPLS6Zx6V2GJIhiL9JnQOcoaCE7WAP8c70nHW5/ogdZMi1pJ3pF8Hc
9MbYJAU0TovjCD8ntH7cFCxC+HTwh8I0xSIea4ipF94IXl7LjKDL9suUgjBNa861SeRuVWq98LRb
w5p2/sFXYmbbtkzAt6nLS/rGloINvRkbKBjV2MpoF69Ndvz9AHna9ldhXepRHpqOlSJai0PtVe6n
3GYrWcZmht50zfvIju1BJoBk8frZlIsFPsNBBv6UB9wl3QE/0mvMIO5oqc5cCCJ2eRsUhP4oxlJ3
v1Ya/OSexSUTAbB2whuMpbrbsuqe9JDIy0iF4u1r6TcOBl5SsCbl3sLwhFu8VZl2DjeENiJD5Eie
rQc3aR1hJnS/UneErX6JdirZb58TXosmSOOfQAKC70WX2U9HcpuKHY+RTyNurQ82p+O6KHfsYaGQ
zVBTm3x1huBoJFo3OC/gmd+S4Zb14tbjGjpxFNPmI9QO3BKf8F7eSnXqDQPoWjAwuwEruePGwDbK
NGcfiV5/mAr1NSQmWUn4gsTZPhZJHeMH+EZBDbkTVpioKTquacIaJy2ibV2xg9X4VrfMd4OqzOsY
o9pmZqXl4229keVFyBm0cOFTqsxrhskFH7o5uEPJkKjLBF/RXFYPYkajuBzR4kL/A2B3Pcbm0ipR
UUVJ7t/PU1LPNwBTmRET7vHEbd0GnODZb8RGAvGhsTZ5jm0CvWmg1hcndVjs/iLOAcf4hnz8WDH7
Pji7v+kQwIuwrKIgV6iRkZfrLogSKBCJPrnHuPkizqTrv5nIwT9JEn2IxxbKdlZsWhGlNmD94P6o
EN9Oi2W/fyUwBvzSKtnU5wLGHFCTsWLHUqBR0hn08R4kEMGEbvRr13NMUOnMOGwAfxduNTSY/DKs
l21YAkEcuUwfFV7VP3K1EpDQvGS0cjg1tiKNuYPjTYLLLJz+d5v2cmbaP+4CdSqkd4sIMUhPJb+s
emu7UW+0Ak4KVdWwpE2Cv2KXdvWhM53BrPZ4gpOLzz/hIM+vMtBhuKXUaHPZ8QF1KlTgdqScAtgl
bUVGbPYNzGlFw9Wm/Gi4/zzNbBkBFgpUYyG4Y1FahuIgiuMUkf2ctU+Su2lbiPVaMc1dLqCX/O2G
UXs4pUQU4/GkGXB3bGvrY3kvrQo3AujdMil7ldAUn6RGrLNFEZZsM9Jkx25Tc4h9FqhjzC3sZufv
OO5wBNvt3/YAEAtpE+Q0zCWeBMSuDRZgA/pUYDRBwJaA64hS3fq5ighXyBV6GZhdyh3hbtu4pDqu
g7Jk/aOAzGm7ylRQkpI9kMl5o5O1RrhQR0sf8HyYCWOhE0SMePSFyMff25zBQCaitWi98hwf95L6
kx0ftmvveGvy8wyy9iAMY8BLWOIsG2KB37L9JEjJLrzbLIkf1Ux+AZmGdHSfesdiomb8aMyjagr+
M48jcL31CC5AVaCfu77MOQPfs4BetOovaG2Ev3iOFc3wxQ8ZJNUkT4FHwiZBUGqE8dsci6AfhTOD
36PKdyIlyJONNoC5gUhzAx8egFXuHvtRXrtP9GhNDcPSc0Dx4ms9fqpmWPfwfql2adTlw0wtWm9b
epQv4exfg1jBU0rqYGtSn37Or70l+wSraAWuf/4q4ccBF6E1l8bc5F++BA08ub6UoK4GqKz/0QVV
sWZM1fe0Lr2RULcXqlh55YKzHJ25U0lt03QFT4qM6Q9AOGXDlxLXAErmkCyiOmsWUbkwZTaw/cml
byWcm2Wly+3unSNfjuL1B4pOEsWHzbrce3nk6hCcYc8meU7bvtSlAV/KuUg6g0WpV5bnqdhSVmga
Y7J2IcDIzVF7gf88M5xN5kIrw5QEpVaGemH/aQeSR+HkdiMd9E+noWi5SDn217bI3l2ABcUbhZUr
b3ldd1hNWdwbQx6InExwd7zcODnwsKg8MPk8zUXprgnYOET9Z9FMYzH23/Cq80K5VLf7w5KT0htp
iiXIwOQ/UgcYvIZ69Qo8ag5NJL0M2rRQmKITrgcqnb8ZPL1V4KQTjVSHvF7vXyptaUT5yzVDaPaT
vE8OTk237L7yJqbSYTSNtttX5hhdnNqzmPOrOZPRxsIYPCYg8ocUxxbeRHEiUScO9E84wieu9Jcd
x5C6H6dcsrN24mYZDhHKMktRF7mAxbO58knmiyhVbUKHaXJZ71Rt6QamRzsfRWedJbMPqZOWGtG4
z01Qs0lneKNzY0KIwBPkiJzvXcqdZ5JdewKmShycCPkbul/x56GcrA7gSCCNOu30v5PbyO8wprMR
tsP+BkZb2E4MIoGowq0vPRdpTrVdw3v6MGuiqe0l9ze+txcPUAiHjVumWxYhvbNo+7rvqtoq8dSR
nPSLyVKTO3CAabnpIuiGly+r4ENIMWhQg31TFg9TJHy4bTkx7pMmaqR0OFpAAjDHxiDc9hG3nlcR
na0o66Yt5zYH/heq335uP19bkLyoN1yAJe9NOipoo3TC23ht1iDeBK6Lj4cbiNp141cJV3dlxKn+
rlhdht2Ohb0xVc6jmJZj947rtixqzK+Gqq7oOLxwDuXyl8ur1ZX3onco8JqQ1PjDAAyCOHUXadGU
kALiU1wLuy8goOkNZnehSxEKdEV5b71x7OUitdLLSDbiAlpGsE7rRu9usfoJb7assyq4dGsGm5g7
BRyt+8RxlhGHpnF9xGxLCVDf28lsXGlZdiJdCihlyimDsO2Brw88KTmHeL4HdgfLdwxf2NZmOTkE
5iYxCWolLDIImPNlfHX9UmBYZm9sMTN8eIQWaHWilTIIjSpr5VEf4OlnBOz+JsUs2yq4eVBr2mNi
Js0dYOpB3SPrRA1IFKyRlaPim3pUXnk7nVPjL5BO4ca1yvmJLC8zKiSXGXdPCir11EayOVbDWm1P
cR6NscopdZCyglSFR7nkSOicOFRM1CtCbPjpTF5L+smvez4MH0EeyTuWXWkQz9CnRdXkg8QWAzzA
BJ/8fenh461cYW5SIEHvwWrFA58wcmqBPCQTLVQMe85XL3ztG3L80J1UDGXi6OVc1ML58TixRKGA
5sfppi6ZZCCWM2hcADYMjttDONDoWfU0oPcFDpICI606pF6U7QkWq7haA87DckJlB2gpIorNgXQ3
WhuvFlobB87/ai2IXVYs+tdUaiF7Bce0Z4/adXrUTxhdEyItFaLWVfGBlJmtQhqAEsB5xJcsoNRr
uU/vlcyVZDHTu5zgQunYwGLunT9IJ3EHwj5+yq3xPhGAd4+G0KMs4CswWO8FBXxfsorGwPjqoH95
i3eui7PS3MZLM2Xd3z8D4f0+29RijjRgF4IrkuOE2Il5UWff3xzZ6HlE0eLMGRIVTWAdIJtUz05V
0ns37L4iVeIOeH9OAGvVpTKge7XBtNAN+52XjB2lh8CuckY13hoel9zrAv+AfEUO0z6sYfvOLawx
ZXrIRIOpPLXXtcla8INIZcHnhJmQvL4Gi844V4BiH1D6VtorN3VVdq8iMlqr1P1O6iDAUOoWSBZV
we3FunP4hb+irCj4RYKxaBDFITunyb2/MG72XjfUiCZQdmc1Hppf1xFo7c0a0YR9PCWZttrekrDU
gENmru8qV99bsojikZ93eAweg1JAPVhUub8gAQAQpLctT13T0+9HwK26bEem+UnLRIZEFe81xC4j
Va/rnC15Y3U00fmj/Z1zf1ZY+8m5hpnWoLeiSBWtLgOEGc1re9NLubk8uANfH/nM1RQL6dN+yONn
gsQ4XBDtUl8HMQwY25C0SsumSpZpiIpcNIg4IE2J+EG16z2L820Ghj392AxiX3z9E1/lxttiPWmp
uhNrR3XQr8NWOgRUwyGVZdIqmamJ6F8vYlFy/nkB1tokX0x5Ks/7XfCddn3EKFHr2bHRP4VrbJau
6dLLYOv9y1kj9sKMws/P2zcqGf6J+PbqS0m0SN1nk6r3duXOhu7auL6CvJ5kiNDyWCKo6UKDkv14
5Np15+lCQzGzui0Oab/Bbe9bC/k4SEeSKH0p5tJ/o24ivGvyK+22DzeV3yBwBpieUGy8NSB3cjf0
ZDs69hx6oV/Xm1h6uaeK5uKHLa7P7tTeXIFyrbIs2VKBB9eXreAyCWx8upVILsIVucxDTzdBzcXd
WstAKcTrlhj38Lgqahj/U1W6ATUCssJix2JM43JoW6q+bCKSmTlB+IXeNCCIiA1OuMKIG31M9nrg
FYZujenmWurmPWlcXQRPhVWCLKJvetmOO4Z9o2+By8YZe2R2IKHAU6kDRVdmEzrqvXQCQxi+YQ6k
3IpYpauYGxR1X8mtO3piFEqSJUVgWwL3BtdNIPIVrDAWTUBaRcRJql064w1yWusXX/wnnfuGhy7n
jOdiVD788pEeMh+q4vjuOoi84NhtdRBxJvLyRjMQGgjdJlgxxBRgvYg8xg4ZaIs1/n7hr5/eNe+x
A3uh/ondWXNUndKfzZZUAVZMpCb2V6ajWK+yj4LqJK0MoltZEvfcSz7AeWnqLlNfBHVvhf+6cWAL
T0CPGV+oHEDrDuJn331dEDDjoIgBPOlYd8KkDCpyhbqbMH5n8UYheoGc8vvKe+QXkiesZRqgCUMF
Q69Q5t7pdFluPUdWbQywRTRQPEj4QBIKElJMuCOll1CH/XxpU9dtsGr8GFPlSeg+IBFcFsLPPT55
U0agoZ9zu5D9qsHRh7uyaP0te1CKSapOWVz1c4vfBZFkbSzpFW4dw1SJzrOPwBGGvaBV1el+1q4i
4fXqUmwzU1nzkFomwhPQR3d33fPrQO7wgfzWFEdHiKsUf/B5mn2h6kskeeJYwXt8jkQpbLXYzQOz
e6p2H/6yaI585mWfxcz4rOl+qPn4P7m52dJ5CMVa+0vfoKHKJUO5x9VIJ9b6EI2xYw25CI0VUyP9
ASkJhK1D+/aoeUjx/pV/xVAQosuKOWpsFCE8tIogOy9QsqLMsMinrS3xs5hzsQqJJ0KpeDmcM6na
F1EP8uFDyYIerfeLJuNtoAYannxHHEKAclK4gfL4o31fv3rP8eegl0xer0MUsVmXzkK+Ux6tF1Vp
bD5K9iXUMY41+T22Epy8xL+XmvwzHjLpoAp0kELB0lZsJb7m4a+RhpNMZjgjGC05UbwGl4dkV34F
s1rBS8chiz1WrRUjxtmavZKzXyueYKQYaKyMuCrHGuJQ0H/1vvRQsk3TMg0oaC3awRWZ0yXEnD/Q
y7BHCjtmrSwSZ+QV0eS1egNGCBMKdSpigcxSuTzwmybkirSYGcJqNP7Zrg+OTDLXkJK6Yw5rbvO/
NjGGz04GFvck32rFyqPuMPPHgEdgMIXAEFDVJ27V36zjf4YgmNwazp/jAC6LF+hbu9rCkVt26D79
QkPYIYuw8ncObVVBcYfcB9wYeSRY9YOd1p3CJO0rxL6ykKpGaNsqIsezmdnLWCH/G5y7lWIn/4sv
Fjp2n50hmjSfWfEl8lwQWBpY+1DjQcwBHRav2YWG9ZikbbOL4MxWLu1/DQVA8zK12dUfGZOPma+R
SetC3ph+IxmTHr8ah4dMqWoctu1i7iXlk6+QoKa24Cn6kxd3l9JGBpqiBktFkb0UDaQE7wctVY+a
eWWKeN/KKjyfHPGJ5dwCd4pn9+8ZYiUynETxLLhP74Ud0zZGhvuBqRwzgCwWX4i2crafQ5CyupLy
4LkUgFjD2llDJNw91ww49M2ga2F2hDphCUtV+2iobCQXftbtzslwiGu+UQUGok/EqHj9hRbsIkiv
/LIN1aoqaJa2B6RNlzO5WgheUYJfoo63sWpMtMPS+kzXlJ9DccJAwFGINbqSHP98EvjMFbMLD150
ZEEcj1jQ2Aqchk/QrxyPgGQo2KMMJ+RqX4VbyBXEJAqn/eRVVj+RuR6z8xsZU77Z72mbtoV2qpn9
WapOjULJ/lYf2Arh22reiRH+DdWqnKjKyQ7VXGFkl8mNN3nMFND67+zpiH+69kn30QcWDxD4uHDq
aVhzs3LjDjhULs/pEVrwyYcJI5cMwivGFJ08KYwWpxUmqgBJqekgXarvn0r5YOHDCLz7+GsE6J5g
fiVIlAjhaPVh7zCYSsx4JgyLHrYhPqouz6ltndMdKIN/1I74rQHZZ41LPVq0VOrEmgU143u0t9y9
ahxPTxsDy6x8b4iliuJdi+p8nHm0X0c5kXIcjlAtuaBoLYsyfMcObqS1lJtGFPeVx9JboFQr1dEv
V9DFi9ULahC8AjEsAFzb9NBM10jhyZLil4tUkX5tT+VJDPBoEIxegvjMFJzCzkAhZda/ZiuPOOzd
/nawmkYpxXvZ/bbCdeLlJrYKGJFSxpODxhx0O47G9pgGsjLZbht4ztee0LqhbMyyDBjasgQlCD+l
1mEULd1BJPa93/lLvJ5jFE9q5h6K/AsFJRmR15cKbGuCQLiTiqeozK4h4GkwRL6Kb+3iJ0nP+0It
PBzvfKX0ZP4sZOs5ro/tS1ozj0nW4m3uoKiNV3kIxhjldfUFDTAaHikrylf0CMg1LwblZU0D2l0U
DkStWaP29+Ih/Gdz0re2I3mMKixLwgQTn3GDUSNnqJZ75HfFnNn5jBzTwZ+sFRxqcPwtFkUryPZW
lveghiz2WaEFRFMXxISW44aMkm+XNjv/6n9QI08a46wDzbS79AS9fdQpxGuPMiAUEhh7sqbZ3svA
0ZblRQ05P7OimkY+rt+5Xn29xrXGtdicvAJSsxNLDx+OHBASmqIbKPj2Bk2p6QX2U7Jjd64/ZODb
Ony+guA2J5kf7hNYeKuBs0cnQ2mwNla5VCzKP03RR7sqc9tPorY6xQbI64MhZ1fRK126K44oD/Y8
OzPO/bpDCjmCAT+sTReDk8pC8kTodjGEQY40UtZXYLN0BZKOQsjopjzFuRo7Jl2817qlcCSHT1Qk
MmFBmP5V2/2i9sYiQ1kwxhcljkTYsGM+Di/HWs+4GsPh6xcGcAZYT+arllzUShVUAYKn/S/TRTAp
SH9uSdt8FLvi0/sHWAaqWH9fpJ4ClKkJYDssEfoWDGAXUjT5YYtq/EBzPQMHcH8rbhqt8FTDc9ZM
G65089E0Bwku2cwK4ylWZOKwZcomUkv3jryvU7wtaqsRxNQUsOvKncdatvh1546n0ZTXO6nmUSS+
2FhT2A0OH23nsEj5A3y8Gz8AmXXdLr8bBzJgbYVYenfqxUtPgIRRZFrchekyVjmElFeyhB8pstqj
5FQsazrjDNUUgc6RCd57DwsHJv1ltFILsyHrAuaT4nMdmUEu75I0owFcVfHpyz5S7HUo3BF4zBYR
Y3V9Nz3aTnTrc0aK+hVzodnr1dGhRK1nXRSzvrZlprnQ6rI9CEhJ2oULmZP6qxLHaMbjU+EFs/Mp
Bj+zb3sorFVJlAXJKlnwGbCvamWt9xxplxvdng04rQVs49x6S2mbAiGwU30SsBWNmIwXD9vd+mI4
awuPACwFtDp1umT844P3nr+riTCMlvGj707RqgF3zWcj6jq/Q3pFsIgdqkI2yPDEB0lKXB5HXWl6
rtXHNzlQGDKmTAIxE1MmObzLaPzsn64n0uouu5nDR1SRnYgcSAgBZng9i0lPx4V0n29OaQyBkcOj
uk8SkFrDLYJc7/ZvrIzmWss1VqMm/1EJ2/sNVbdDgtL9/7069eUzW6jB81QQYPAOqd2twZCb855p
NpfgWssKlwdkcBRQnQPyV1jWsU+wBLOGDq7+fQs4+32wBaL582koa6yrsm2trC3gtOhaISpnxFbN
xSHbB+5sxJezPnstolgWWiNLoMiZk/RUSqHMr/tu+UD/zQLVm3jNCUa2KkqchglG2UXfY8Wfi+Ua
73YhrxW/1WqlxZwoHzHHfq2VTMFOI3ZSOeqr/LduN/4anj6P4SLj2vbknVgQqyCZbrlh96ULiEEx
yQ3J/WiTMs2WpMUzKRC216JCt+Ge/1bv7rooF4YvH+4AVneQFulIpTL5ndbB2cUQmDAIBB7+W0dA
iXyvLyd5NFKhpA+tbRS8an6wjrwoVw9o27wwGx+z/Y6P5ML932K98w5vDJ7MqrdhUrNJDwCwRiaH
Srdd4jrIlENejo/nJKTbzqmsHM8pYRaD76odf7zbF79afIy2HUVKcewKPjIGANtAeCgvdS4TdKBT
A6cdbt9ae7cBrzihYFwyfBqCdBOBGoxCZGB/ddFVHPGUe+cqk9W/BIWv9HZ+7WtnvDcvrFxbBv95
JPZ5e0q2JJVySpUiYNtVTpy4IhBqIz24Zyr9ParBq+YY1zedIeD1g+xa1wO9AB9pcaiwSrS+0nMo
dEEzYUcky43/qLqmJpmnhCf50JSCNyYu39orQ78LoAWdloc0nJyMacwkc8uwHtuG57FCcrz3HL+v
vYC5EXS//kvtJjsXKi+Wapb/p6N6YsV/5y4pp1vXmfEkxA+AsTfRdL1w+gveSQNlkeB1wEi+R19i
ua29iMVDVUp9GYuDvVTuO3qZ5plT2tB6o6AJvKInk3DLf29pe4tqJ7sDZyFDP63ONfx4/gKBM+s+
JlH9hGMUUNhcf7fY8DQ0AFE1g7vBqqdvbUprForL+JiVvhMRAjA2YdAxq4L0UKEFKey0MEnnBPiP
4eS0YrRGIbfuAVkmP5XmG1JXRtrHdLkbvOwnXgGeTzxx64G9m8vZ7/OuXviW2xcC03yl5PB4twA1
BmQqhW9lmeZI9b8Kr8S0rTBytHfDCh+R1Y4j9XSTJVqQWEoUwKf2WkCXvQeLcjEshdplRwm1/zFl
JLIkugl2HhWX7nt21orzWIfPSmDLCq2LcwFn/LOQID+XuH6HZivJu2gqjcoRRTbH/OhVdnvWHF4Y
ZnRoC1g9kO0Ys9A0kdrIhoMK/uvHa7oXoDJStjrzTd2Pn1BtWvUsfwWDX60mZa+HWObHsEdTQpqa
i1N35iZPQkM4NDx0eF/+ShtqgAC64sdRkFhZ4u3PLXaC3vpq0ObAsK0F70KfxLIjeM6zeiAz9bQx
Ci6uhFgST5Q2vukI5WSJRkK9fiGKmm5MBNL9xsnQQ3QHNc/fXpl/cTOP/75asjwQaUtq+FLqiscj
v0NCf41lVbdsH1WAMD38gGY6udLb+OgpyEB/Nje4ypfUqfco/b7fOdf54T+XBYH/rsGlI3Y297dO
iAHa59f58UBOONkWSjEXQOeCsSGetBzVjqM7x1DHdSfZR1m4gZ2gCffr13hOvnlnOME0loPNWSVE
YPpahE41DhhhcTDrJxw+iaxXBEqPpEaVFPzZEMwt/OsGv5zDAvazX8a5OaaJLs7hGHA3FTP+D9DJ
WG7gMeLN6yspk5sje3DZoXVurCmZlvYa4XDxUVbwDPRNDIiYQJvZDON6aLrbMCy3vseGNDA9q8tK
trdIydJCMoczuXF0p2y29jA1DqvL+tESTS4Xrzra/AdFJCJMkNPVTH/xxzCVOB2Q99wCkzTfqVWM
msMGOl+UqkxxUc2sUzKjNNh4Z2slvVtm+7v8MiBEXUfNsSMNr8scRKc7LLI7Nu0+oNMdKFthEblC
Kw4T1yG/eO5MC6rVRfR++9IDx1QF6ciDEpiIceqUmnsJ0nAMtya3Gx065a8uF3tE9J+9cn1YDCsZ
HaFI5tM7kJI2axVU0BQQWj/u6LY+MA7wpRzwgJWbzA8+lF9h4Bkd3X2V0i4m7I0MWMvVQFg1E0rM
OWx5Hlfci8khWRAlkxtPWG/ULJrsIdiDQ1EB5nU19DRIJ2KKRkHYlhTiGID6/diCVNBe7xTanlU6
Q+DIZgt9G0ysOqzJDOMsrYJz3BNy6cUGXDa/J/3oVpzyBV4A0Bv4mENRbkAWp3Wx2l+TyCElZ1vD
qLjOuOYPHq2T/f5T+0C9q+RSmTViBJh1HoVz5V6rHv6xBuVFpA7P56dXkef7NEzYa074hikrITOy
8TcVZ0j5TjUbvOqBfHVSRp8FrccoRA/tgXhstz4hyZLP5cX+cwbUinDQekEvVivfi0mYef84caSy
9l4xGGpG/rAGSWjnZ04Ch7lzN0jAf8hGlqFXWOVnrjfZETU72hU6dVXTWzIXwpp2Ld8aXoqbd7kw
1Op0sTc+19ecbzaOYQnyQf5fC0IkSO6VSc8saKe4KyorTrVwdT6OP1zI7yMevIS9l4TGf5fEFREB
w9I4oNtcjWr9DEc9fzQ6HB4Iceu47sOAgWVzheRItB5R36m7pFaua3Y3Ze8AiP4kIUxrExXNPSM4
d9uxA1FvAbI9FfI3jOxwSaeRLQYrxQNNZlkoocA25p2y3g50+gwV+ALEo3ZSaoXeqzwPCDPwZbAJ
JrDKd63f0fiaP+6RZgwqBHchXMEhfVmJz0dCxn+jXp4Qm/OuFWl7xJWU9md1FZ1CDx6MoNAz/NDz
x6N/6kNaX8bZj4+4BFwtj/bM3oEGkoAdlZG/5DtlVEncrFLw5ZfqnZtofT872beKI4C0f7L9Cksg
O+FCWrPn66XrLaW6717jznu3Dd8gYF8cf/KOry6DvW0oubLrEosGPSc6Liq+77UKnSBunC5RuYDI
ozHsWmh+Mj5yh1+s/lsCRdh8r3YdVg8SaevUFgnm2SrdjZBEOIwpURaQWYR9E1BGtW/z5wGw8LuB
/J2bC8EAiyrDlV06cWWW98T4bJAYWNTwuwbjf5PQAkS4r+jHLTBkFlw4nXe/LelSML6ag3kXj2Mj
DkcRwdkjfHXf+GbW8yMqvWHwFgeioAPADuypAtAWFt4tmZM/1lBLWJJPmOtpMMRd7eIiH5xvmHtB
BIa4B78LCaHd7CIaGfEbVP7vLOLonW9Hgig5h9gTL1lYEtdrWR+9nhOESMcEtyaFhmAYpirH7pi4
FyjI3vnA8mzE0ajHfuSqNYyM4fRjzU0cU00C3jdzN+QaWuldJolS8O1k/g81sBLDfq1JeCW8PFp0
UpRca5cIqDhP2PbfmoMjAQJw+uFFWfTHfiFr63CVyEJrRZtiun6DbNH/FsQ89GAoGFEHksAACL4g
MFRLTowSoT5ZmvWLejkMqDxPbMzgWdy40Q+gVqE0r3tJfA1v1ahgH0CAYXkBRtcSnTAhkQqXqMF7
xrMvQABA5uxquWxOKNdTpG6L3A5h2ZjMGXahTfj9aljCdTZwMXDdk+SQpskOXgpFWC8KumZYLfCA
yQQH5PX4WnKqzQIFdrzVLWwu2cJIn4AAVFlnbxKY4VfhtybrdC+DkDXKrHR9S6xCvtdPS6acHY1x
ccsqEgApxbyZrQ5u7fmpOapwKSF7XU1DU0hnRhnaqOSN4BaY5qDcBrk/e8MxNwbgEXahENlvhpaP
wmHFYzw5HV3vtX4+PpozfzovdFusWHzO8tgNP2wngRdck88PU3acDYGsMsbOa1YAI+Rx0qvoedg/
MRFrOP6nXg4s3gBxyP8Rl3Q6We+oLNPd/dRL3KwPfL0aaqJo3nvRLKKcqCXEGoLhpDynnN1ZL+nv
DJm5+Cr7afTlaPTGE7ztEw3lahWlS9e9SLFcgCXs69DgDfDVsp/d/d20l887Bb7Xgjorf/jvI4KQ
I+YedqQQDgkCeazIQL18zaXPpf0CFI9WPj2udbk7Karn9qUkP/3hdRsNb26S/U0tjPcVY4uWYYAS
3oOyTGKvselReY4hyRa7PLVILnERy0CrQb6rGw0TXLP5nlm/HK7otu+hpTxVJAFLItx81HTzX1Ht
/lriWfhhcDn00+SQZ+ta1whA4SvF9Xr53wg8zR2jAnXwq0ROX8TGY9zaxn/8WfBrnvGJfsrUQexB
x3PUJj4fchIwWhdiMT4Z9V6FPxEwlxdcvx9LnnDs8WRu7Zq8pn856zxCYqFHmRcFj/tifbUezhc5
KAivCQ2MYmlZzxZvLu/IpDbUiDPoKUe0uBjXJHWS8CrnJSrQ94GE4ps6kteUkg5IuSXIbzrrwst8
PyXIqcR1qObTi7puMZ4cIJ+Ju2RlbfXd/EZE6hIBiM7n629a7A+a5zjOLlmaadz15cnxhUYWrJHV
iTGdnKgj9K2I9cVJmixQzvscEoRsJropgjTkC13Ko0W0O5lAgh+aHe9GKnPNyaw+EYt9A0M8pavy
cDFXfGWQi+AHPQtVuJTNkDIqSfCeirjDfj6VOsRV5Of7zq6bgawSlt6b8v86Z5RwtTX8hwORhiPg
SfZeupptliHqsOdskAAjGhyNLo+v+0fbKgTHxMSfG0mUnr3MW3otgzv6Itj6qq0UvTzaXJK8MDn0
hrNWc5BiKqLaIITamQjM46Zu4UJiULBfpThx8ZKReAwDs2pLOViFyL8RLk8hlvgeb6yTbI4qE8BZ
Z9Yeixl16S+RMpJcaNgiC1ryDAqC9tb8YCHFo9o2MVPkfejNA3pEoZChxpDV5+TPdfIYPdYwezcQ
3+H7pE0vgtK+HQ5TWnhoE6nEhQDK1G5UJT4QbbPeUaZ7M6/rbaXiZWW/9unW2STGTSalXe2KhalB
l6ox/BN78RxY0eFA74BfkeL9kZ6A9/A0s1DqLNQRWXsmSScfb5W1vMM3Z4FZ2LEQNxMTGdsfO7+f
PH0kQ9eqxfarOtt705AckYB1z6TMtgRgHz1fkNmWvKZ0lBtVZSi46Jpf00tTXVA+YgjQDWxZKYaH
tB0arVmxIdRHEHQAHiUedlkkgmpDPv066HmZ7KfWbErg5ehhaagHAAizCytR69eYbLDkV8CmEDvh
NkAJ802HS+0Fz9TvNq+WMeqjf+C4vuNDmTixQyRcTXrPkpi25ePsK6rDNkySq5ScjfnztVpXESPX
57UNgPwJgMej6oXwKfAmXM3IrVCrrIhtvIsiwgRWw+EDZaUHZcLGxDjaLEbK987klgY0MErxVhqt
P1XD1Vbt+3zQ1JM+J3WaIg1g4B6IMKm0dxf0lDcW9zVKMrnyM/KDSLi5/wCbC/OCwZGXUGPqP+oH
rOmBD3ymyF+EgInfBfRazqFlbjiPPpkAFHZ5urJ7nfWCyXXRprSfBzGN+eukHxZfUt2HrTzcvXo3
LbGydDzjP+udej8ffWFvzKOPJ6dzUcA4WbuDbZzD7DV4MQiMnVTSQyKPU/h+Cgu99XpiKMjLl4X9
7n5GzXIwh2V13YTR1Gujgod4uIf4lDvzSRyVkRsNJKtM/H3r34PJAeVDHEYLF9+XoGBf5mkl45UM
TvPgXawXoWVI/1krvCZmlu23fZ4sXN0bIOKiJEi+nrglcT48gticHvJ9LmTQ9QBshpLWCyBgmV3l
lL4cUE8iY2V7/KahCwoiHqIG6krceC1rLi4K08i7srWUUrojXoHPZ5ju5oSEGTjLRAP6P8vIyNlC
lDJo5Aziki1hAERu8GcJNPw3vFiBRPK1W63ZFHaSiy2eHyozHgRZVM7dsfHaz+gPdLtf99FqQU8J
A2RR8JCtOfo9/3psZObz+WbvKlk4KFwG16YY1Rdam3lKV8QcsTpcrl0t6mvLY0GobCoWPhVLPfv9
xzukrxlIoB3rcD52/ickwSnKRvhPkw9XcRhjGw7yMF9XbE/iEv5BPUjZBAqxEHkLCLkAErwrLRUK
iqeuKdTZ/7iHt+k7DEqPT0orzevKiuuuujeQJgYlo1bRo6DuFurdy6e/Ren9Ra5W0a8nR8PvHkEP
jxfQulgpEyvmYFyYbL2YYzJ8+VMJql7U3fwoHnd3h1uOGJXWZDpY2rS7rEqmlTrK4COo6W65sC7o
DN/rVkCLgjazfkZ9RZdvAXoVrgLbmrNy66C1Ak/yCfPXDND/dEEt2f35zi9edrZgL+0FLgHttAHv
o61f4c+Ocpju2IiSZelbY8BE+q95/fGPgJtznOYzKzlD/33zfkzsl1lty7Q8FVA3rn4J2mTsoEVb
wpbSDjDDpKnetIZ88eMr8pteVUeoaPKZDX/m04kadlpOcUyrSUGBFmbmT4c2qPDJS+1P9O+B6Qkh
r/rDzE5Pq4WJdn7xAw5XZ7ibba9YMuh3Neo2kxLKz1b1HQ2OMvFuUGBEcH+9rGyz/zTD29NtQ2Hu
O4MDrbNECtOXb3le0hEClmMjNSS50k+yaohefslVabMmeCzI5/ipqjD02d3styzFLqoQEKrdY+Qp
SysibArqQEd1mEcBe8Va9NSrTwc/UwrVxQOS2Gx/lhE5PTrVBprTVDnik51SPRFijhptN/lAqobp
UOWVqR+VlzpQrqRO0eqoB50p6jJBTNDDRwTBOswAsJ2oZJz47Z6P7lB1zZmoB3eiNTjwoJv07xCq
anEwVwGZmxhp0zK3JNtld4FVGPN5relu6ZFtfvts2v4UTnu2veFqfBtqoBGqKcR3nlQYP6OvavE0
8kz8CYAnofHqwQqrRKO51s+nYJjPzSvbd7Z1oq5NOsXF0+sNOvOhYGy/teoeqq23vnSqDDpvyhsu
hSoHk5F6CXjG+xJJBL1w6aoXCD/kl9dNUYwNIo+m5z0dnHWuoLzjcOEBDwONwpplrbu7JruSxpDe
M+aqNNxpgftTv+3eTmYhAgXirDksq7THlzKqBY4Y/CfiVnwRQ5NdN0BZgTo5YZl5c8nyeNzezl+o
1NDJ/Nwgmy6rvmSKyEcTGOYpFkyuV1qN0t7ZX7H6STFMGApGm6lk9BbnGGE0PpJqrsJj2iZSFylL
Kn4W7JPpEb2uRrpMEZJW/l0mMeTkHVBR3kRgQPQs/qN/BYHkmCClpQIYqklD188gxzyupbDog33D
w/8sdLXX/Z02mS+Kiai9lDuS/59ny1EI9HnSGeDjvyl2zDyS9xPsDWL3ZzTDiLiFW+0kpGCmKXtI
bRA1cQ+SwXjWMTLsFcr3EWVvbaUtSn9zagU8sYNqj2H3R8+/2LvAKgvrNHmnAi7GAx4oHPPHSHf4
vKdzOXGzEOgHsvIVeLE23vSJfWgnxLcX0vqGOor3I6CV7SPLkskK4CCKqF4qVxuo4nxDeU5yj2PT
SgETPJlcOhntliXf0o2yg2DzMtamgdtxmI9DMi1LNFTpSfe8uRHgy6ps+mo8AXXwyl9qQdYvLNZr
ueTNic/eRLKLSwQlyjheFm2jeRNYkJewXlgIQXTfr2z14jjf9s8UPdB5kWwFthiFtND0/tA3NhH+
t74h3GHspaV7S6XOzL7sZ1/Pe20YEKTN9yS0NAlalmPBmqj2h6/QHmckRxni+6VtZ6kj4/tdsusV
QsDWWJSCW9ld233mW3PoKMDoDQ7aGPfU3BMy/OKR+/txcRK3GB35k/HXZ4eRpmiqC9scLjxGo5K1
NIOYZuRjscfulLZ47JAsPzdgIwgFQfBIbEOgNZQ5i0pFq44mJrAJ7om+JtVlnOpoj0zi6mZgevKv
AYJ0Xx1nyC3EkV8fmt2U1KEA8m8bJHif6sFJh6Ep9UaLkcSuhY4DbnWEikPnmgbduALvGLH9P+Wm
2f0b19EuTOU9oEhRdC/SgJaNKEj7/74WL1wfRKUDZDJqmPywi6tyXRpuCUWxj3gqynzC52UI4EeI
SAOWtfZvOS+zyjl23WQDyyCLHsDY+5+CwKiyegzfVhRtNLpvAh4K4/sj+rq08dNypJ7Di7vI3+rG
dzRho5A28ZMaPPPzOip8Qlhe3g9BopdlYLermEVka098la1pYcZnIhZOvVtRC1sTGM4xA57kx9Tf
sq465O+r4sfrjMZSxgpm2vXRLomN3jBOmEw6qdgZxwxQW4zdtHezokM3Ug2euTv4trjrPS/NtncV
u/R3EFKbBwyABRw/0XAG3nN5FbHSREp85Zpk5JLsB59vcorNsDsuD/6MYupLJ5byURQYZq6IkFeL
0Jz3/9Yp9UjInetwIal9sFCiFsWXb3mNBqNfSFWTt0qS5PxB4Oey7f7+gMQ3gnxuVQfsQTVsO1uM
aUtjOICehI0G/ZFL2m0nzvZJJ4Q8Bt+qWi+yohoIWxz1tnURrQNzfK/Ox8woCx1CCXrbgtNsvKb8
GMEjw/bxNjUjGqe9N95pLdmjvagBNLexuaw8kOoXrTcMCXv+EpvmN789lo0CkP/Zg9SnnH6Z9kPh
cOVuc4tpBTUTuogoqTy5peY/NXsYouyT928snDU0Q6qmWnKbOZfYZXuHq0WxwA0UTsf0ezvdNgFR
Cb3L6Aeu908vrKNDiXuSml0C6gOBh58qlhZsF8ZKngdhDED2XpcjE+AHEh+xaGaTJadh2gnTN9QC
o4ZIgJHPdLbOe+AS0bomvDiuqUbFZUGPFkrG6AUK16DeOP0nD3JnEKsAPrMEVV+vW0goN8HREEFL
w+G9GYa8hITqoBS6+e7QdC5d2r04f2saCC9agLgQJVQDxcIU4oazDzFFxt1QxWS+/Gt/Z9G2o2LA
pQ4hESd+yrOp/WEzIRvTwhe1WjzkxNuExbKPo8tengm5DoW8rSQzXzTaD9WYp8LZlQ/L6OyO4KXh
i4KIQ1QaZ1antOa3lc1dMyhcEAsAtIgXznY1ilR/S/lvsuuw2FW72mxhqpoi/Zm9LBqQ7FnI+ibS
gVNisucackU/a3IagOZANHtLCFGYK3ifKNk/A4flUGoBheBDcSnMksYNZ27v/bHGYMRV08TqrlEX
VYAlfWXICrsQ5VOassUeiCHx6KYR4tasYsmV0Z5zIAhyJUaVT02jwWQg3w8DRBvz5uT72a2+IYol
aGybMwbGTkoJEC+TVYzfAg4QINrvj2OT9r1WpsV1CWkOA+zD+Juo58rRolezG8vPandv66IwnlSB
T/t1TFc/EzHmuwVuCD9MsxAns1r0y393xmRQ6TAvbx5+GkBWYnFhqgk510u7swrmR7YOSsQtLqQj
NxR9MFG27pCvihe59fnX0FUZlgbBedgkxI0nAxhvD1mHIpI3RKjEMTKMCSalJovuk/0JClLwpxHJ
f4pSEu5I+/VFEEdgDXwJvXZyFsUVbNdOFfp/JlxWI2LFiM1ZB+2MBi+6hdrpEAdFBFMbcG0Wuxlb
8x0ESGawxPVIM7bI0sOMjd4N47c8ae/bGXWSzXUDOHOREOMcgyIP6C06MLkwEVBohAhYwSIR/n9W
JcXQe02V+2+bzZ+YsVsz/w1HJVSwl+cIFo+aMR9J/Czadyjhk9tMeiEQgAeHaS97FPy7r6SGORda
yBQh+cmPnLAl5BRBeTFoxoOnnNsCpNzKri0dLc/b0s0hqog4b1YYaWF9HoP/eKsJOOdoxET30P/w
+m6L55N2Nzx/yC0SFh/qrGrUJlpPWu5QKvvPe5aTXt8h1jz0n3FGB1KBca2WRuWtw4elDVO0rVjT
eZ3EOZ8+PbQdj3bKe+LwwY4fU8iDk66CKIcqZFczhmi78109q63Pjd9Hs6bVI8a1ToU3OHyowON1
CvNkteZBwJC64vtd8ihHxSzImTnXRXb7lAVoT0wqegFk1WFQyMyzh99dzLiO7/1s2ZlMA9TVrINg
xjSkFAMC+baHejuMeLU/Iv238YDC4U5QNak9ksVtU7/cVpP2pNsJ5aYY1gickHabf8KEhgTYfUP9
4vCFMojPV7QfG5zTMCa44uHAoj4eIylYx61Jhpwo/su8qu1bZMRKfzJ1iQJIKF3DxwzhTRgO3ddV
gdTFIGuOcJ37nFy2PnGZfOEwwoW+vSpTMeW1ilH0SwnweASJOuQHI6plmr7dYyR4QtntG/uyngWS
xoxsUtwH+FZZQaUvet4Fbq4rr3LPqIDAhtJnpsSrk549U7T/N7B0UDboUCPkzOn7CigwO+hiWsY/
Kjoe/B2/I4bIrFVe1jxjLCpSCqZoVJkny76RXOWeBYOtzy5OwXqrr5/sHsp9SmJUC7F2tiVf1rzd
fAH1aPxJIT0JC4o+nnarNf4WPep0MkrjlBGDz5TCIBunVKRa7BDEnaPzE8qM5yNYF3uCrmzg6VK2
yiBfVNaHYTLyh0hC2KTFOy7358Ti2+Phj47AaadMPnItSn6RTDZ3OMx9qqgV7rrtGwBGy4Fcz8oX
jCXX8jq22IK6LmNaf/6BQhOvNq0u8L0G07gg6xp8oPV24YBfkTW4CHcCorp/SCt9SeMIT6UApQOX
ilyTZoz3AGruIR37g/e18D8oZj5HhuNI0sSwchf90MPrP6l6SmrpF4P13ZPylhgIAyflVvq4uafD
it5+kTUPZhF4tuBXdKid8smOezb6kTn2eoq7fpqO8kDPx1s6N3xJD7U+8wwr4ijb4DOW5r3XBJxl
LZ0H9krH+wEZKhxnphEaO3gi6YUfq1DrpXAXa8HZLvjS4wRdZ9fTmpy4cNgFM+obva4cBXYo1FCk
yQNEhn12HtjZlkcna1ThnvA6tcYU0S621zTzbKPsDoYp07QFzTQdsz00qPwZWqCJjhiuBm0Dt+Wp
lFkDrt+dMirP6cFyiOjp1mSVM9BGLnhVjS/K/w8JwxfWWjB0cS+9FGliyO2xBKuUuaWJJajYu4tt
PpWxeC6+OcGD2xCWtdqpOqCCJcbVrfNs5dJaXYIex7Gm8FoImDpTMhuuX2AFD4p2P0PM7cSC260u
dOdzNcMNlY7uHgPVykixwUrrUPDljumZgbnAs+s1DE8beRZAB8o9erA8Lz2ziHXYSgYDnBre8vTw
IuseJiv+Fv3KvjeJPl8LfCTMFvO2m9SimlNrhb5ywvHd+ej4lsbtpp9mXXrc6KVFbo9Zdyz5JyfK
z6493wZTf1D0oRY5SnmFeequbhIIZ+opjYAepDKkpJGL4prdn/9Xioy/GhYGKHwhRgjaWEpCSPqn
+KqLQlMWGNlbY5mi+ixznptvS6FpP1T3eX9J9gfyLtBmz3ByB+ztf9tNn0oOQeOJz8Swl5hsFKqT
iGffmeErw/R2vaN0w5CNdsTWBO79tbJzZHEHyc9tBTD3dMV8dU2bfgIncQmvMxM5mmfnWPUERAFh
smL5OVVbYRkueJ1VdOaNxSkuwyCh0zD9Sce7V5Tl3Ekc9CWSK6Q5QAcZVWbutATnmIknla0unfBs
vePUPlw3fl/PrDwK3wjYuCFLWyPgx3HsPQJe0y8/5xHpULyeOFJujndPQnNLaPZ2H6hrFfzuuj8/
IOqWtX0AVqRpCvKhgjGNNm6o2TToXPiMp/vZtmE/bDYr0eamqdsn4wnNuPE+0g77xu3LjKeO09oa
GHQoy5cObNKaRESarCZ16QIKiZMX0CJcgQKsh6zYYBXwBD4TJABFLinQP0lFfE828rnatmbRl2qN
Hj9mhFwrsMmGvmpH450DZXQOvvPYo+vnwWV1UiAsWI9d8Z2qQ99eXNc78HlmwOY+XcwWp7uy4+7J
5Yl89M3dvrfbtCRrfmPsWd0TuA8Nk33S7WCohL8Izxtg3XNxiy4z6+jqqz39GFX9vk3iAtgcH0Cq
m8pzT38yfXRI2xxchEownPyrmYHeLiNyLH+Xkcg4mOZhjs2r8IpoZncX8ZOJUj15G8BbH8+bWnx8
+1XaFlC1PKsT7m809A/TfVFWIrt+/tFI/jY7cCBSp9SjSQb+yFjgsmIlMsWfgV3h78hi/pi8ETSX
SEtv30KfNvaO8soLmXMj37EfB772aNRoSr0qmGPlyjaGDHzwe97a/tqdaSuuSjDBMjrdwqvrPJya
S0fR+kQJQaI5aH8KKubohU2ig6WtYM3LY23ePkKdDlw8xl+jGcay6WVR0adJQWgFHT9yLnEKqusW
jGW7l62LM95kkG/tRcnyiTO9/5n6HyrhSx0YXuF3R1C6RzF3MiepAXvHvbg3xXbbMhr5emRaQZoY
rEmROlbYr2CM5vwHih7GTIA1z8DpfHo9lt0b4uDoNNdxlOxZihwrAS3+uojGDvSRDEmOSdw5ssPy
YPcSTDYaTJPBJkXTUSsEVdkaV2lAaZ3VT49GbP9Jr7c1GX6Q72KH0FU2JBWA4PIDJq7WDeawg7Jp
tAbf4outqzjlHe9kNnqccqLVh8dCxFJHO9CnP1KHVOO+YJ8rCrBGOc4zu5xtnUrNHbddAA9sX2GI
XuBNAwyetdVo7RH3MDBjT8tNTZsxgv43iCuWzTBU1HhJ+sZBLNxrzoRoTXcdXctVyEtvbWhnEawI
xFtfK0kxKCKMXWC6h6760GyRHfOIqOItaixuah07+8pXi7n25l2/GG/G9H4x/tgAKlxWxxMfoWhQ
g7SNHHFLx+8K1u9OdDjhCUtfof9MKsz8YGLUra+jARgTnq/tPuKjXwL+NTx9w0DzTMO2Mh+TcCeR
iD4y3/a8CyI+w3VGm1S3Fk1Qc8g0Bq3Pwo3IpiddUnN0uR+44fipR0QBeI1IAgFPFw0nIHlVFkw1
2SLnThM9JUK6s6m9NwFM/SwJrSdI1yp0VOyzJr6iw3lhlOAw7Up+SzO6FeQqtiKyiWYLTpQN0Jby
DpkiQkhudLUyHc70tc22Ef5x1DZJQkJ5zBaIVcp7R2UnIEs/DI54qNZrgXRa2pn2+YKbU8sBKayt
ZRNKnV5d7Lt6hhjDJ4L1xLH7Cd0MFbMynts+zQeszb4GZQPAnV3qcK4jUzWvDazPhguoWJX9A0Aw
YnMAhj5CO3eGrmR5xkWXuyJZULqkROFB3E1o+0CaagQ62yvu8M8io4HxatdSulGdA/Kvc5H+1vdy
Wc+PjYHGWDDm6le0XtPyp5CVWXCsV4Q4604UqN6ZyfDnE2g9jS5KGQvZUcxtMRs9qr5DjT1kh0V1
vJ8V6/djNfbQRCcLVw4dtIVzSQwgeg/1Ek603Amx2pG1taKCEQz4/dQfaOa50+VX29GvdTDBfiqI
OU6mY9SoZ+3z2M4cMmuEkskF8TpaBlOflJEeprTPFRuhvZF6B/W0+xEWZQCYY6c8+R5obAlBrKtm
PZzB5/EENPe0549GxDjIttmdmZvDp9tk2xGpPNGITrPunJQZzR86MtgqEIzBkeJOh6J/hcnYNKtS
Dh/Q44txSvo7JkFRPqXngXBnYQoAJibM4xi+tUwe/6uzPWk++l66H19359OgWYlX0rt7uHTXtjOx
8UCWiRL5tIGvg9tykQOIgFRYRq4GaucJANMKhhcHtucg9SAlm4WM0WMnbpe2kLG+4emHPsqCPPTU
0WwLqUoKY8kXAucIIJMZQPg2o0E8LkAC7WQamehboaV/UrB68iL+mHafFTz/xFmcfoKQJ8ciF19r
v6fjyJQ16JjAjJQKU+AFFsaj1nH33GjXmbU82znMihYfw0IDzob3Ol5Q4izBrU5B6Lf5WQlOxVXN
iq/nO8HiC/InDdqSI7Gi9WiHc30o1t6HtJ/Nc7J8OpOQKVF8SxeQnoBwp2WSkrG1HnaVL6Uu97RW
LgWtfZr0o3uLYwuyWWdo618Yr7rzL0hCoiabDVhnkI91hBZU0pU6sclAL3/3Sg4sM5ucbxDPnhMg
DDnE32WpAyNnFdhwuUdv3AsZo1YO3/mDJQ8VIrCfoGXyc89lpfgt1wu8XjyJlSziJXqQAE7b1XVH
P3bNlKcafuMaT72YWiHXeCf6J+XCvZH77cjJgxZ3ATZKJh+V4HgYga45jsJnc0qxLq6sOiqsuH1i
gX2O2EBAsH9ODCtkbLc0x8sXLytQJsj9GwLYCS8gaSXTYKLuTRRFKHw8StVYoWm5b4cFfmOyiU/B
m1r6SlED8VdLT9/8JzPC+yJQH1zwWG5IlUssAAaUQaPUkz6MX9skawz01btPqZCtTCSeZBF6ynx9
OqbVSj4odO8H2sSbznWljwJT00bcs2r3ZfbcTp2oUSlyBQIpMAzZKmq+7m28tx8zs7J3c0K+YZNN
3AleLNoScx6lDXBDInjni2K7wSlm3Z71J9P4LkIuUPdCcfWllM5+l1JRboIaAa/FGbiWVidMeDqN
DQHsc0c2OuBEuouxY/E0cXUrzr7T3Pwq3ek/oCWn8X1NKem+SP7AKpHQPtposhGAVs4mlFFWz0y2
dmZUjtE1V7I4tbBK1CSF46u+4dqNE9WDDTDAvzl+sTB7zCd545UaU4xcjeVJDMr40HKvhO8wnsta
i0X94+7sWdMMK/uutbpLww6OGU9Cl3sTOwijIyj7Rlr7y0QcQOT1CVsKwICLj3V0pERMV+q+D1mV
aUtHAF2QSNYQIAsb8uvsAZklfgEG6eMc3BThNyIwQwzLJUArNIX6IjFb9p7sBsI2FUW6aNIZkueo
QCOzgsKejzmEZfAONj0r6n8lNPaCL2Fy+6TZz56SqYcPvOiuCxSLLcpQ9gvM3vG3zQiAn2H7NrHK
FMw3ahdZZUL+PX5SyHtVPblrLDbIvnC65LQDMbtqXs6g9hFkjwVA0wHRCNx7xtzIuZpzIosxe5ov
VLJfj9M8Jq91DOLpo/NwM76ksaQUWjvgzGzHLAgX8cSn507DuGDNN+v2E63fQtwitwvHQdGfhhN9
4Ls192ITDoC9viPTQCubpKfiggS2csDC4WGJR3eMdzqKbM0DOVLU1yBlO2FRxTxQodL0Nhs2gJwy
90sXzuOVvbGvLoYDRlrdBnP+dDnzd/wbFqlcDU+it2xb+/A+9RD5TmspIGbGM8XQoLGHwE7RWkjo
K7/Iij4s3H3OhMg4ikJcj4qN5ENFakQvThMv9F7FrLmg1oI1+IlXgBjkz7Zi1SB+TWmBQCWh1UAt
2KbWsOLKtX2UJW6KA31ykCAVmQkgabNoidLAn1fSy+iY3feoGWCtaqpnP39/5pFQ+WaLhiwMBtaG
1UCr17C2/g2EqpkHb1sdo/y97VlJCabtc+7gTZDBmtcdmu+jSf0tvmRiw0TYr7lUzV5bLDohAbAe
hJciFmyt6LLOO+d6qgD+NqKelE7zRLxS81nKSLTJOFYLpZvXkKYnFJ/svlBOVGMgc9f6IrT1PASX
pt13BZOS6CUmqnrKQqDPOaeXS6N9lx4A52rGugZ6fU1Y47L8fR8AEWtbFIH0vNlxa/uVyGAOWFxg
H74bxUmL3A+eorUJ0osPLYafH0lxYJaQamYlsV2Ymhr6W0eJQt4AgW+TEj2+BmJm+OMpo4UnL7vB
WsmkzRS8YZIVT7iTNBX5BFL7ONO37yqurTzIv4diR3zP+ynn9PQoai8oknMI+UjrPcKbWQnVoH4z
A3udlyT6oG3JWoVTAml2DMw3dpAqPJYspwo/SEyPxTWZuI2Xc3Ue4qKpK/hCe/LwetKZc4usToo6
cAA9x3wGjuWF5TPsif6txe6/IUeYatpfMvbfg7oQ4WW6oyD9bU0kYt7fTeDzhiLVCyxSWqQXZXW+
Ns3q/rrR3bpeO0AHmXl3NHN6KCYZ+nbJl2qEuA+grvBJCB80ZWw1sMGsXvR/6340/4ask1zqhsvx
TJGJ0qFdAwLuRRNie2qr+CJoOPfOT7zRYGUMZ4FavKzX3OcVND4lA8xlSDx7wH0te48Mjc2cG5+U
+lEdikp7FvIFH0jhniPISS603pWNCdB6Yfal9VxAfpFKf1K7XLVJhW17FSR5FEYK5sb8IKMMCVRu
4how0/A2J11J7B71609/xPXbHm4oBzwnQ5BwJiFtYBrMmlxe+2zk5HYtNNH+LwPGEDeB5/yx0tEW
EWD3xMHmlIK94YRFaM1aH/PblSCwGp58ZVsXjZ1pwzrVVsAlqxf6rUA2XZsUNIEvzGTP/nDbqLRp
8V8A4S/Uc8DtBdHOfhZUriinnbPlaMzjR/rOqG46VWS5YkF+B0dumHphM+E3XGpETvxohNTVLmnx
PFb8wAOOtLnhQYYtilDj47FkfdTfaCdFNec23RtWaqe++Ex2fPTeWURlc6XXND0abbkma43LCsXR
1QNjYo312VanQyDL6nPP90Aq1MYMmBokvUFrckjz/N5aX1mRNkLu1rIW4iyTjo6xMfg7mP3FL8LY
JZq3TgmXCz1SVNRZUyozSF1wsvci7WowYb8K9ePnXzXpSbS78EyCeI+/h5/grOt5qToiaQedTHrT
3/ofNeWHa1eNDNPogMP2olPj4Mr/fiY2Poe9dlHmVwpajQw86vf36vk4llEcVtCxi3UD+TyUgpev
xoNK2VaBJem/KHbMZLuMSjJKbmFwWYAdh7R5C/Pqfzn1EPoS1u2AMQT2nf+J+sGFtwJfWNqYVLXz
pDTu0fMu4zZw+8YFYui98aAr0bHRbkySQv8DlEpyUnfNtzLaPNGwJdmvyJxLifgeWHMaItVFDxfb
I2XuyDzb4esfoJUiPtfdSK2A7sHMN3zldUWtNJcA1fFjaY4nxJr0eYoiYAY5Op/TJsthzFMdKyEM
Q1XS8K8M6wrf8gSZ6k5PzpL29FTex78jvmpdHZBX0j8xF55Zf2XkAILMG71gl6El7vkxDVg7P7b+
KAxN9t9GmL2RETsvDLWmiyTfzIcH2aVodMv+2E3uQTXr5AA63kKH7CsFPzkOY/JxE2pO9O1WD6xX
RZbSgG7ciR7ANNd5JKeZt5ZmajesCWlID193sNMJJO2Cw9kzXqVodDO2xNQK+b9Ludeo1Ifh2cfl
9U7QzNcVUoV1givSiqg+1KeN2MkTQ36SL+PffU5C91OlS7c8+AIvT11yv3XbghgbzWsQQA/kDkYb
Cl1fZ5y/7EZa0Numlxi03gNO67f8epkrHW4HSOX0OWH5Vwzodhnha+kvc8TGOd/4pzAsPeQ7wBV5
3G6P/ucmx9AHeMv8AkG3J0N3j+PNNDslwsV1UvPYqoBRUvq3YfCRx1qR83+KRt/y1w6adQ7gHUNE
GpKbrPEHWbwaizqNvEpOlw3/U8X7uJmT4rEaa0bNAI4Z+d5HiIbwEWyr5ORrMzvVcbiNsKsxEUsL
EcwmjGshmZGHWiuwq4a4gkYYNsMpBAacIDLL2PGc143NkkfR8rPVNf9pMGP+lCF0FdXY8Pz1Nwxc
7+72TLuiHkQBXW9KT7k33q5TN2W+SsRh0+oTjfgzy6qTfIKyMCPr6GiJ3a4S6yV0F53+MOyz3X8P
rdDAMc7Sp2+My6ZyZSu8vkac86V0j1gNFSHl3Ht6zqM94bZ/vMSOXqFDDe3NBSNU1zYG/v+A3Ncr
Sn13M8u6uENLcvRXVRTevLBE7EkXpCPkEU6MC69DkU6L/31/aUHpjsNOM5FCpOqXdeXm72+nE7sb
JY13PQzaN7AtcEgWa8gsrySPo2oe6RL1yC3YpgnEQyNjej2+vjqYxSGYu1BZBYt7BYE5rswJFhRC
8Dij0Pfes668wCBldXFC/eM75hJUefCQhTgn+tpXdS0/qIMmOGAZgHYQ1HcGdzhl22ahQwJH2ZBF
caCkERM2byKL4q4oTiQz+yrQHoOhqb9CBwqWh/FU5xK5hKiXmiWPP/5yd+D1vhBoaBFQT/6DhoIo
b17bT7Qq9U5Qpo6VsLiB2gc6ohJrXN0i39lIQUZlwYcm0rrUXaVP8FXyS9HWzU4i7v6KJ0UjK4Yg
XfR1OAclQrh0eqXMYiUlEupk4k8EHDFF9x5QByUcayz3onCkrTECl37PI/Sm5IFcYRcgsMPpslgs
kXPeadXCIeQXtAxGkgpjIB/AP/lM88fD1dFqVOeGHyYnC3iUEBGZy8YPYOmiNC937r/JIRdqp1au
QST6zRunSX9FvLU3itqkaTZuvhQitGTSP/kWmFEGlXZe2dUcXQdQNBoZWifQ+MuuR91sTyPnKfm6
KlZShsqBDFW75tB0UOECzrovNwhdcTuRvRF3VlKBxgwbFVXt59AAWO+Pfnk/uE8et1ghfaYo3Gmu
J7xB7R0lpujV0DbHI8MDYfdy8SzzDShQvNvRzupq1EUtK/ttHSew9/P3FGru+tTwjZIOtkLzGtM9
aQKLRY1W70bmqW45W2nTI7LCgEIY49/SjW4uLjnN+xcOQgPsPaLe8/Avl8G5uFhFeq5gmtPlA5Tr
3BjhUXzKOADE16+AcDqZZehBR+cyKkivNaQwgelQy1CbsMZuhBIVs3qiqoCAvr6VswCkaDZG8rSQ
oB3R952NpGwS5QA3/Hm/nHZp4QRb4knMdODRzBsMbGWYRVuT3YENwY1TqQvj1bnnxqNsblnoXDOZ
p1nv/OWkm562SZj9Mw8cS8YszlrvZ7GotcglbGXbjpL6owE1yf3q01IRgr16ZnB1mU/fxZn73Sz7
5HLfxO75ScLGJdaubXHlG2SySsRiIBUnqU0XqRPBtEhUAuMTeNOlQ09+I3nsgg72x7O39LkExH7n
LyBiKx7bXOOdPaS5Bp11q2AvjeqdBCqCbaCzP50ZbPIl5v55loZLabKG/676/XkyMx4bvKY9ZofD
RF37ovZGl9aERl1WmrjoaWeeW2ug/Z8mDiNRvkBGyQQp6WHQLIAbR53sqHQCVHYlbDWE6bAI2t45
dxgCb8T7zlWuCHVQ7RrXmKPZ0RHonZsNf2GFtJMA2ByyjGv21KPt8TeS21pOHp9jS3DjT7szxv6+
fpwAUOJco42tg7ml/OKq8BVwmHWJZzkgzRsNYgVtOrV0BDR+B/i/B+pskQqyh1sNT1yO6MDXP0GA
qn3g9/88MaDHcj++bP1JdV+b6wLGmHeGRt7RWIuHUwadkUxHPCja7WJ0gju5KXY0p5oTfAlptV/+
HJeffo3bVIdkbmZYL47bzbqm3UbUYy213Jr4canuwT/pzGpBWgatiZFww+WtWrLQeUxK6q7VaEPf
DEjp8/Bt/4onTVQ2JalUAqwB4eugiCpP4fXRy7gA5+ua+4ra0rkZINP7VNbMRmAvGaywisyOqyC4
+uuF5DHvOqTOD7ar0Hc77ueXIoa3zIkQZr2q/sNDk8WvptdtCdH6WIugJIji6c82dy/UNoXY8qjR
mcsZ5KuJPv9iQHcEzIsk5AS2bFz1Wyk7pyugOBBXUyzcCKzlWhEMJW+M4YgcpQcTrab/shLy1TtN
gJCbTep/qNO4h9SX29pXSZHmLmoGiCJ301HGFx3OxXGi8M5G/QJ6tjReMsGrBPiArEPywR0J0kkk
cGdiUaoFT2RWGONTva8R8jtXj/jQWYzTpH8Jj73OWrInFAC5TqDe1Y9FXkIU7eYadUWlaXIUt+kA
qrZL9e4WmcISW+I6P6zg7EsHJF12orF8oebhWb5dlDGtqHRqEUUxuh44H8g9bM1B5dxTtdXnJMbG
i8nOJl7ay0unGEqYP9z1lOtK99O+1ipb5Ko7w2z+8jYE1TwJvEZ5pvd54PWRzghaCWtzsewA3QaT
hXnwrGL4ZAwo5rFcPmxxnh5lny5XqjOpkGaxQGPhoMK3kyvhHcpstRTD0pWTBc0pfAuwr2poqAS1
Yz8IKJhB1hkFgTG18LV8pTUc7kebg0ACNSSZ+qXU1IqQNW5LkLVRzQcQNDT1MgLoFmQKFYm8FMMv
/gJ99VxRQPLLGhc9apI1Yh/fKKCyhZ0soaEQ50nutcAQXWRY+ck2YGf8sbiFc76YfxYFD2SiTTmJ
UKN6K3OHSMKES7HXUogODm5LmSKnoIbHcvFnoO4E9yO8cg8NP31OUzJxH4LancCvZAGFboYS62C0
hh9RhnNriVj4It2aYe8bmN/E4hSSXAoy3qsCJkFqX49OTaptdQy0h2zfV4MGYaVVO2v9/L2yFr1H
cTZbNEb2ffIKQKhJ4crtJSwwpfie6HlQvreoA34BgoWm2oqEW2+hRLLN79jOpFfyGHcOikSt3Ii3
5rLZIBl8bUseByC6Z931a3LC8pjHuIC+wSMbaAzNgCtkTvgXXa085QTC2UcjtgGxei49RuUh78h4
QDGSWlDg0L6C+0PRLrEVPxhpVMbrMQr8HtNSHgXpJtl6chZZ7xi7j8vnpuFysNzPy06+d3qpUzC8
r0ZRSWjr3s0kFuw+RVHWbxUMG9EE45Kk0xHtMTdvE+uEmkk/2l4TTX1R67wuU843oH7mqavJ1cWI
30DV050rv9FrdmoIslDmm0N34VAbgdi98LydiHInriiucZNsYxD2H1uZi4oZvQ4vxrm9wXANkL9X
QR/PYu4vV4Yqhjjp9GyJtyxdpeg8HYr5vYAy9sRfdW5D/MHBngALlJTg/3a7DI7cvPsn+2WKJYzY
9J/62aWtCtmWtD48brmZMW3hHgrB30D/ebuFsU/bpsgywH0zlzjxAdA4LFNDag76ZAKgDAPOVEXz
Kf5wG3DBB8+Y74Au8uad81uy93bdCuECgP/WLTaojWtOqPsQxpCKIpfvHg1UYMaDXgVXXvTkKmhu
2A7puy/zDzi6d1seGQCPg8LNRCXa+mZ58JDJfNX7PHD2lmsolasyWgaqc18pJI3bvQqwxWYY52ZH
HDd7+q5KRTqOO1iZuMfxjLm7XUaI2oToCLZODdaPO5RmkbJwuVgcCBoX1uyvEK2P6SygFKFlZOzR
XLQMGlY6aXKhhB8Vf+e0EZK7DeMWU0/kSeRmwoUxRvKimtky/tNUYl+RzVzeD578H+mfvYGX2DkU
ZbiQyk5x6zykpj+CW4kXvpKx2ZsikPrGfyBWNOZWajevcEEElDlXO7LcmB60HeSHY8GqnG/6he9g
AEKFM7Bsf0/T7kIsuTopsslLEnksCzMy6LtK5mr2Q4kEDVOwWVlcpqaHNFb/xnKRXh38MWybRG7l
4oRKRmjavx5MxCDTlB04c0DimzqzSV923vM8yecRQo6kgL7FlhjnY7hp+rbDkKw1/vfZzVv1Gocp
y7ttPvyTojhv5Dg9vE+B5ro1WeoM+3i0xt4eCxf7Kt/m9//4jeT8eziei1l5NQ2LP6mtBnTFPnLo
F+wxRmcF2Fk3Ov/sIt4Uo1lUIQjZsSafPgIDochgpn0v3Yj2yVQT3UvkHtk7e3LxbdmGGVPId4sq
5rmtTzoR1ovc+Sc35u4WsEZt5uF0tYq015nHNuL7ivwtkVIKVhApHC4IA7g+OKb5C/tNINe5Ma3X
7zb3QB0LuZTA+kamkmtPWnw5tjhvsUh7R8LoVOj/TeUg4ZH58c0wKUZh6GGQW+u80iIY7/5elRkh
2QGxdZBhGhiKJxKKNt1eGnT0AL4AT7GhjVr7JzqOaDETCTWSAEiy7aGEt8NV/WnzSA89pGwFHmsc
vz0Sfa4dToBP7pG9p1GvahMWks1bvdBExWSG8gkUapkVpiIvK+Mf8fL57KQDJVERaxgwouPi5Oqo
HhQI6cZV57jxEqTTH9EV0+aqEzj9IMRh64NzJeh4RoBi+grvZMx6V7TSVsE1Eg9LvLN1oZIFrMTK
5DUfk/EK5PrOTroHEFhCRlU9R2U3edRIdz2jlacjeRMG97h/3cwMHYndilpsZ2E0QX4OhzNtW9gr
dOmNWX7s0YREPGB1GdFDtegiu/lUqIrGPwZ0RnRP8qzgAheUX/eQRBDCNK/UYK+1B+ii+7FTfIlr
7emrRWSuRywsyJsnq9/LZ9rraEJbh/0E9OXWNMw8Fio4cs/hFNhr+dza0EQ1vIPuA8CNBIz+Ci0J
emq1rPOpC/W9yTYH/YFDyX1wQxuT6wCImiDQpGpmlpSWM5ZBUB5CQLjEWDc3bXf6E7FNDxx62iOj
x698DtaT2cCnJLgCATcLLf/r6T7r6+FUra1UbQn3yFaUUrsfGJjMHwJ781i1KAUyiJn0SYp2mIjL
3I8PcTk4kNUbga+eI4Qg7Qussh1LwzErlLEyvWICMwB/qkt3bfTxq6RaOSfpIWI2Jrp8sES0cS2r
h/9ijwtwWC7XryXWg+NTTR8Doxptv2WZgQppGVkw7TxgHkQvUHCEXQx7k8WYpSEfIxA3CX/QwUUz
5lp4bDTyqEaQgCf/A1IEhm55OthAlUNH2OzdrFQ3NyoPCexQIzi27LNej6WtTC+7oV3l7fOP1ipp
fp9tS8jYBcbI7EdlkKnhClKct29y/W98zcbdG75LRAjjakZV0mGdyVJ3r0ZO3wdewgZmnr1F3yob
YSCsuhsm9Vh/g9LuKLRGeYVdc66tz07OftgiutP0V0hGTQy5Rwb8otG3g64dJGIFpSz3m2Jcrw/K
BjWnx00tTKN6a5SX+/O0FlN3rtycg50jENbbW+TaVacGgXZkqGs2XQEnBDggZiL+d2YKoMzISRDm
+o3q8kjKrLScIGS2+MF/jAUKXCwAYLvlHr6QMVG2gy7gDsYnhtvO7Osksbvz5Un+eiDPs+9jZI36
EF+mlniPRvtWSgsibWYyLQwc4whpx7GEvVDGIwOrqjITspnm52VvkAqWpV7JGbkV5YrFntARY60l
dKx/wqkEmR2QcEMi1/TdyEjCBXboqLCuU5EBUCqygQn4t18HQW9uD+oO7P1u0LUa6c/EMtRDVxOS
YIfXFZBy5+LtcNPNmOlzCOC7PkffQK4dP5M8u3ZGDdCWH5Reo7JgzTWosrGf430JK1xBecaS4Mbi
BVaRTfVYixOQfjCWZArqiOQ78ElSmkB0K0UXtRmXVzvsT8X9jkP7NX3wsenW5Mh/fs4mzHg3NLSd
AbYpMw7bBT9MJ6s93NrzSdYM+p6p+xZngVt9HX2oDd0ioTJfZlJaQUG4mQIARE4Mtav5aW86VOyX
yzalVAT9xmSjKVKhzTqnnheFZdutqHmlpbDSb8JoygFTtrcpdIev9G4eAIE7sz1bk/XPfyaprGKH
rSfjqoaSIeGowaPmYOtnxiHqdFL6tPj8dp+Rongb5lt1JqewEI3VSGYI+wVAgA8R6cGZoU4LH0Sr
CU49wJxRP7Xz8sWfBJsZIAzz0gtYzKuuaf31JJoJIHjHLLgItIJaRNyR82iChUpVy4xuqMqq+899
gh7Mhkh4nVK0g0sBUH8Go6ot0TLU3A2BaMnhDLJECE85b+qIVi4z56bTDwzUd2w3POLlyC5d10PU
cM6xW10YtrS1IhzL/RAy3OSE0OgA318kab8uj+pC84lN7Psq9adbE7S48sWI1ClkL4//URIpcydv
cwc7xXck1rJCDjtxrycqggMpOWvIUprNk0Za9l2DVvggqOXym3QW+LNO5F99fFgcNLFdHQ4rkihs
wt1w0fa+RbkD9Gj+C42jNFV781Vyficpd10QGUiPpbRRqz/lZ61GwM57xoExFirzobx7pktLPk5K
jUD2JV4Wu+i06znKPjyl2jjlw1YEqUDfCkmBF7D4VhdyMykboA779qP+6aH6t93ZEyyVl0OxiXrw
qWDbRRHZ01hsskN+x7pLyZTwa9D7di/S52DO/pW665TGhVjHfxYUPAkkzVxziUOHeJXEhIjTAq5m
g3nAdToB35q6dAquk9feMUlLczpmDdN3O1+Yi8BUGPzEccGTErt7xYS0mKIlCzU2LBAowCbMf6Jj
SYF6XJQ0CTmq5P6PvS2IA/Ofuw2QyxVlaGyTt1lhMEoCKrS45e19jP95gyV3vFKs5Uv9kZlrQTXa
mf23HieG6yqql9S9nCkakzASGgsCb+hAb/g7NI/YDd9BkBKrRyD1g9K0xFBgS3rJihhdiQZirLpb
xElb4Paphgx30VIzZriftAZoc6ZuGiOS+Gr0rloaIpW+DiE7ilE195WD9qP52E0oYpFs4KYF6Ol2
jTOG2B1mk7ewNM35tMkIcG23quhSCwP2N4vF3BIAmN3TJ+Q0SFqgcCqZgcd7gUIWuZT+7TyxjyjI
UDv7Xb4RIAJ0e+tTr1dwYKei0F9nvCrE5BzcnqCJ3zgJQy0QJ08EjUdYdT0YNc1jb+Pw4M9lqOIc
TAvZmfV2LJRJjCVydW6yH6ybRhUmcM/fyjqEomguUPUm/vSrMX0WTq2l8qIzMvXpwRdpUElc+Jw3
hEFhNsLaJR5HVxSydHpMbEjrFoQu+giBryiONua5qa0i2xzF4loWwC1J6h4dlORZzRT4mGcKSpaC
Ym1eg3i89YRge3jZ5mqhfOgpEWESVzV1BwMP4LZPjVpuUJOzjyjRne91a8wCZhwmH6ZIL6XFgeUe
oJ0MJQrJpjKbZjDrOHQBK7L/Tz2ldM2XR2y8DsCupa165jhL93Ye0B2kU4jr25MEfH1BJc5SIDcs
v5whnYI2kPOQl60g36MlSpXgraeN8VPgWv666PhhHC1HffeBGHBbofzvXOUc3dNPBD+Tq6DjPz5i
l6K3M9iGV5Z3oXr+oigPO3gF8PnuW5QV83qm8HtbTcsE6I2C/uxT9uI7mroxfk5MwulgbL+9Pt9i
BW15c+mq6rv3RDei/C36xY86hQYT3Y3ZcoMjg39/Crtpiq75ZyJl6u9hTWfzU31F0/z+2iWYiMfE
sxMq4NRa8+0vh6mEl+xZO+HdLV9mKSiPWvdepI1pznUykxxSnOVfkoRmWWggR1PXARB/GyTD81mu
XWelsx9a2iRzBIjdr3FfK3ZXN8L+31TNKN+Wzfpk/bOyLzRz2J0CXxsJ2Immf1qCpKo0YL+o5kO/
u2zKnGSODudv0Y4Z0Z9jlPcI++Obn6wlUKauY6nCNYTvBjyvnektaH1TRmOVfUJ9/1sm4eTOke0m
DgSH5a5I0hy2EiG4qTHjxuRDz7gMvajU6t/7muE1HfCMj8dATmTraZtTljx8pY6apGC0NwUdlkXe
8I0ihWZ8ZTEyDVCKtB68ASyZix6GoRa1w+vFc59yUWOlL4sjHfTiUhvszE3vWnrd/J52BbUHWqXh
WvThJXsokXTttmQcgfBTdOQEkQ2yqCGstyRhZuD7JL38kfmqRM+Q9+1viSYb18mNLXnkFNsMDFlL
HaBGIzfGEPVtk/ZOC9we/hPtM8jHxGkMmHgDatK4uUFH5aJ1yjR9bhsn7cCbDhG3VUHjCe/t9jXd
09FKQqGSaq4bkPFLy1tKjC+HFyqTIkfhG0llp5RlFBG5kFc4E5MgdU5XlAv6hIvm9Eqf2UXfnC7i
VvycmugRPLwSTIL4jxn7qAsULLXIxbf8xGE1u/aRWamSb3Ks087HgY1csJ7AVF7J2MRkYqLwa1xT
sMMHUUrihUqmnQpkc8i6Px9iu/mo4VcSM3ej178quyzhXI4CsdwKxxoPoLgjrUuElqi6Z3Wnffjh
QkQXIVRBy0SC1jBEs6vTQMKoKfsvcKj3hn2O2n0tzolRcO7n95ZqHXAKTNfaJKU1xJsTdPW3QMPk
7WaXQY4z6fE7fc8Vhs/Qb3VLZBGHP8LIvkq4+ZoWeXqYhSo6jLRz1Zekxe8tgX2Jlmin+ZLR2BCH
cbpS7NDXSNKU+euwkscjH8InMRspzIUOPgmwv3h++S5EsRpSlgvhj7gZ7kxEB6ovRP4XztnbTW7E
RVxwGPqmOzoZIZfmi5nq/ZwMPEpZlIObP0OuvzyToWI7RzYtmziE5BlOXS0F9MGK5fagsDfyKBW5
QJahFr0plE2/04n2HoNhmclxfxbV3MYnu0Xx9fa2sFgR0zCNdVwCDx0sGkJMW9V8BPNYUXu+kvDO
+vZOJkQuN6D2SVb5dsbPcbWOD5B/DJRowxlU8WLaeeTSBLUsbAnffzPTRa+FQQ6bueR2Rd1siwUV
g/spu0jXRwoPX9gXJX/Pqw6WiUd5ffZIm0iLrxifaeb8oMm8r5D8szedPdpQv8igmusDUtz9v7a7
N+n8ANjry2wE2IBI+y6NjB0ZkbJwfnwD7Vc32Q6W2qRv/L6fK37FAHZdcbDc8405EXzj4MF/PON3
8MhaUnFMSCwk8W3CXeFLHxgUXBpKuuLMDAfOmWdSMH8cWe7efMsr2wjoGSbT2nbiBlNPrmmeFp+U
XBGdtwr68/lbjt3QK+gDzY+5NiafmNb5I3ylQ1QWlBmNV+owxu2wBSUKCtnU4WwIGdpZdxYPyyTY
tf7dC8euscKPcIOlxQ/fT9iCnvIl2fS7KYFqJe96lMlANI9u9iKrQfjR58rS3+mMJRLcfjR+V/t3
b51aVUVQwFXhC6Kd8YM3UHuEqQTHWz0dGMfTiGdqEYDZO4WkKKWllONAfvXw/8csDeF3NyF55A2h
VFPiRpzJ/E7szzcJysUTTuJLUAs1/LsyUpI2Ws2/mPvbYLFqpaMGSnrPQzbf5CBJS2zt0HFdgi7O
gSm7fd7VL7EtzHMLWTbfbDa9recsLhtK+RnIopXkIoqd0zps4ElYU4xLn0HzAjTx3WXyHEQYxTTW
vw/8shsnLitG2/BirYoW3MyQdUoNqtYk889KenR57vhOw44vjDmbsdddZf8bRAqfeDHqJIWu9cKu
NUbjk8TnEo0oTs4+Pix6rchtYz5uUwQGA6NCy6HYaEyTHZZ2bFMwHcB1zDhsEPO+lMKf5WCGQvup
nalUdnIhsAoW6GlzRN0r/Dy8e9DSAizquKH/T6MYULSz1j51kuHofQ7rcO9m9g0+ohroplR59SHc
WURFWcXjC46KDG5Te7SdX4KkoHMjCe2T7VZywz4/slp8z0vOAlpUp9bOOOnIuMi3gOlkaiEFfJY9
uCfCvleZaWVnzVqLrlMtrF7ZlpmfYKMHPX8BC8nXuKmzYUBP9ABPoXrTuhn04I8cwJFC/JVhevBr
VLr72vx+m9emeSZq0gX9q9e0MaJpAX94kIXl3aV7SCaBaxkl3BLpneSilJWWvcR0V0IzhsyxtHlj
qicNWM16xkIYS1Afd/gI4Bvr/RByaZbu0VA1WBDMhUJn3F6cFnEJwz9ivBBUvAgWzmqW5DpH6oiT
AxUBhN52JWMkwr+TBUzvPa3STe4bsE6e/s4DzqSlFo4Ibk6zsRdJEa9IhX8Ftmt4tnHoOLt/Ey/d
bFC4o7YUvtRLSdQMsvqwhEQoPhU9uIk40HC5RwkQvgciHMIuNK4et9sc0lQ1OTIqwWeDMcFLDdtD
P8bV5RpoPekgpi7v7gvS1SKt0RIrlz48bxNhXChcvaBi5s+XVCr8KDUF3dWWc0Ku1SUoJYaklMRJ
WMYJSHRePtbhiOugO0gah9YxbCd2P5a4Y/TdKelYstUtu1AHEsqc2putjLJC44Ntiv0qLbFyrVnD
CMS5G9KzaodyhC0IElr5qwhGF7gK9IpyqpYhvhHZeFfiPaGJRlsasEvsyAxJqfpHmVdN+kSbXFuM
BTcaSyHG7/oSVimlk0jjYOu7dWLZsPP2L3nxqSOBQHSENajQRW8x4EiXhEP3N9cpvBf4f8fOoakF
6XeoVCQaYZrF2oU4BAPffU9K4y1Fqpie3ehD95J235tpN4DShC3rMowSTriGqID/ivTiNgzoik5Z
pB65hntcp6cZAR5tKQgJTHvALnXPDjONqLFzN6dwrcMMpnCW/ffZ3Q/W1S2Rx3PzoLZGra69fKmL
91de+5ux77cLUc8I3VY9rqITNClr71TobqW1HdsasFflutGLvqT7YcS3z+QyswwCxISQHARxDiry
Qbte0fbJ9Lnoyn9i/lvduoyZNEI0ptP7JwpcfSDD9BGx3OT8fYc0tx1D7G8PgTLNIS0USJM9XP/C
tOHushiSqiifwYFOLMW0oNJd8c0SJIf7O/G1NV8hOiQDGYuz9FglJa3l6W2oo/GgeXmNaMo2qzyC
tPnX8dxvI5uC8YB5qPOytSqte3vLiZCtmEK7uDqyDzDX5WXKLsDsPIziG04nWfibsm0N+2C4dcNK
tgfd/6xCZpY3eWB3YqRWz/N5+PAJD6EMcnoSy5ASX5ecqY0aW32bxtFeQ070xHugGPcmCsGb+FRw
AjQWf3HzRW9DwqfT1fdLRFd1mpPlWr4WxyDsNbgoLbJtAHJy/51T337ewo1Kqxmy6KGxfq/xT8Z8
NkxQAfIPDZJVxXMdLgZhYofhbIBGDrL9gnQT8GL0lvQXjN4UtdH7QihkNd/FdORbgLCJB4r+kfbd
WQFdlFmI9HghDbLdVsw7N6zoymXDfnV8lDAQCSiakCks6tC9hufSIM8/A4FjwvOghK1b4/Uw5j62
p2q7OuzEmPG1wZSrm8XvnWoxvy8bgWmws4Tn/KCHKzsED9PGqVEPI+sXSYVdiGIY9rypEkVNYh0T
TsBbQ9Lxj3E3LKjaCoFJVs+d3KKdngiPs8GRzizS17CR7PH928RTqaogFoMZA9xrLUjXZH+KZcN1
37FoBRbeoG2Q3FUMW6t82f4EMme2LXKEbxIMhocJvOUeZ6u8K5Xho/gAIJeHRtb3PtOWqOurHBzz
vuXZ74Ey8P/sboHxlxXLwRyGGi1ZHvPD9rnnqiYTpLoVI4jcOcxOUkHxqjW2UMX537UPaG4PhGrP
3ZraNe3cDPAN2EWHHE+BfUccg/KinMBUNwy/ZnAfEPziFppvKyMez3++zTC1agQiPeWVIPxsdgR9
KwALe7gKmx+YhH9tOyzEMeLgwjC3rwKMDhktX8jo6ufNcavSSe3rGwyS6M3Zg4u7LgeMM6SzcukA
8lFaQlyJPm5JCPSLE9/Ngw+/aaH7SsvglVuAgpokEVvDrwKhkMV5ZICNwg6IviQAfMdXnqB5TIJE
gycWVKmRmZIwS30At321ftM76q7Nzy0xWhu9KojBxVLpgBSEee+ZEbXAHuZ+q3RNSdo6HmyhI9xg
KwebxYAY5/rjUDkj5xUhAnxiGx7/rzClFdxLfL72/F9U/2DGZQD57eWVtI/x4P+xfmFXHCO+YjxU
86k+dIwhycfIvaHDCnvpSg79dRHgRNBe8eO0CNf2quMnTIo32xBDFiwJ+YiGxF4r5FrwoEf3IpL1
MFIRyZSR5yiSRL/jFXqC5hg1HNkihW1N6oPGeXz8gTWqKMjoAHWMowhF6INLq+I5+NG7p7MnnHg1
Os/G7vQGP7SZ9+XBtAO7yOd5skVpID2BIGwLJrezoWadghdbOvRcB2gAc+F/dz8fklGYIvXEpfRw
3gPQVQYVNvbL7QpY92NFvjgid7L0/p0vzK1oW+FJd/RtY3jeaCBNCzJXst6kEvE2AZASfnA1O4XW
zz3dI5g1+ddVHfSDWD8+mHbZ0vgbQtq120XsF16OmuLctNo3e0MuaJaToSQeeCYZx2WQOD8n6zpI
aaASyTcmCw864ftN1o+z8zWKR2qeCym33Zozjy5RNcS6lerb04t/hEyaIoUu93V+gl1wLPXvVUKJ
mSWtb/IG1Nl9rMLjS15OYY1/0X6NOi2JnTK2A2IsnjTlvU8wwKNClbuZuOw1NDlFyGOkYcHYLEIk
SIxd4BHE2cblAmlKeSGZORr6qtffEaOVYRSulyNp7OB256Dg26Z2Z4iVVQ3cFqDAWjXCQ1poypXI
vZJavuxvVsPUpFGOlNI7NtZNHAjSSGtKOCzNod/LXdWIgFIM/EMVIWI8NxvlLCtQRl08Y+UKZdwg
+2hVAiVcOPxnKd+VAm3Zc2eX7MdKu1RgcUH5ANo9VEjPsPn0n1hnaNRV+ePENBzoHDDFwVb911vL
xh8f4d/tkREWTo2YH8XUdtvD8Y/Oo+mQuVt865p+R0icq+yPqC8xMKNl8JQBzat4k+q01Ch1bJHO
SxtnSVAmRG4bki5g4cupdpjrTsHvWuGNIbEa7JnQ4B4oyp76mDM+guOzDVYmCoCSWEkben2a5O/h
pCTmoB5WeYRhddh574E0U+M0UQ0uOly9QcVnygL3ui2Ccj3WMn6SzLn1wWSh83Hl5JLkDmbj61sW
/fSctd29xYacVcZ9y0qKliwlRhPCQBKS0hRzPxN7b6pPaBcj5BWudHP7aGOrwSTO9SEe00Wq98yb
/9rLnFzfrxEu+cYBRkS1nly6+EZSmuVR6op6+kvY89oYyspJ0DwmWYlpiyk2DBKKn5vZg89dKpgh
Yas3UZwRj2DjxrD/cf7nzwV3S6polkAUF8ZKxVBN8EivZeClXcjBekzfssoq9QGnqlHlSney8n2E
uXPZh7JWjUQJZPMR8V9K0FNtfFC/UkxLo1zOR6CeQvogndXMTM6atEVLyV28K6oZT2IJiWePCmcD
R+B1lBpRiNeEIvYByrY402QNhFABebfUKiuQjcaTVApXJrfC7rFOtHh28VVwRfg2NK6+4OpnxhqL
kTukKfafaGDLWdPoHYDZY2Axmet1rRD4+9ElpniXYrSrl/A70Np5fZCo62j4C3MLyCl3YVCArF6+
cR7EXMWoaKQmHgnc7jrk31Mw+MYV3VU3VXzcxxVmD73Vd0iwyabWoBYOhfBJthrJ0/OQP8EQDGfj
4QFjz7xRPLoognM15KjMCeK6Sn2L/J6qDQWH/SQIF/te/H4LOQruexn3y94+AM4axOsrrLoa+aP2
D7mI6fzxuUeYVbV0FMQP3J/yeSXiunlxT/hDneB+oJy7fPMaMDqZwhWNOQAWI81VZOgpH6bNL4mC
yLuZVCSDcYe2LrzDNyKISqf08SriKg1FnoeuSAg+HbNwz3KSTD+plgp37QpVEZj6G3q5knApcuq1
A8zlk8OKzhZ6COgWWNZKWB1Gft6fv7wnmtuunudEZnPMjwJx4iZLSnNtY6nGqkxay9iEHuq/blUt
I3DYQnFxInGpeBJIRQqQM+Bf2+OZdBigfN9/fLXpB0/np9Rs7AQly4ogke5HMH4MyajPJC94RaH5
MwmpryVvyL6RqpF3YYq3ArqJB/Z098LmCMDJx/8r+GKhwdPbziv5W4EjobI61eeUBwMrTHMDCbHe
kzhMwc/E07T26pniAQVXUs4Vq4rDcpcMUPMhbNN6z8CzHvPt6KZj8ecotRYLkt0yngRxKYUURy67
5qB0TUBoScmUcP9m7ljslEUV+ugnQWheULJYK8tBnc9KvGNmrNW09s45EYqreb1lUGXoJV2FL/mk
KH8rYpUoRwS/pFxZp0eRWLGJauYiocXLViG80gy58C+RgZ29i5LM9fnBNQhpsBIPIWVa/HU1vNAK
LYa9moEpiN6B2w8blfUQqrbNChedabyBb0dRxLKQIwLYDd993s7q+mD0dE32GOidfapxCy9JKfgW
hTmgRUeaUBoO/ZVtDPwY0Qnm06sziHaJGAucH5Aikbvi2pApgh5ocm+oaNbkHynxZQ/NxzQp3dqM
0rTUC/yORHBXiws+v/GPdgoVejzxnNWFE2jCo9DHf6wTXerwGtX1mi/OF1FanaBRKLDO6RLz6vCd
GA0ulEA1+NDCQc/9RPU9pApNtwMdwZti+b/P4oy1Ngqt3iRd5tN0uWgDouss5gelurFfesXpVRyB
+iSJfnod/FE1JDk5yZhk05YchRdUoDovIhNuq4CyFzY1Oj1Uy3yDONB6ztLCZHRUDIBdNrtIDzRZ
uL0L31u930WhNMfTJaYt6ittCF3bmqAUNzB8BXKVH4A8Z7RjVjSDvR/dbKBbIMAYsSVbjFpQT781
iJWu1mEAi4NR/Az9t7fXJhxyiZZl3e4XzQh8CXDLPl2puzbQl+GGoVC/eYqqRH8IcNKGfDgLcpl1
qidU2mOffm/cY65FMN6rn00+ydgcNmNPA3zwvGW2g2sm5WLS4AviTdvzQ26yTrxgKfMwNiOaJCal
1hteHIRh0HxalaEBZMmtWDWjmdgBkeBHOZRvDI/3bqcNiOeLozEFwU6lyKu8nYQ8y1S/xLpLGF/u
2l20NOzloTLcT/cTpLBTCavRC6fVf0IRKaZ2wSEhs1CaDLTM57JUKwtEvHcNPbvOKyurL20OqF/0
wlmNNhSzQ4CteaYE5byp/l0UR3rYmooZWYSV+57qq60AK6C7BAH8unEPNEhtD/GDa4PM3BFjMrqH
fCebw81b/AeYl88Y+6eYVMfHNoHc7BZAksVtx3kz4q1dIFeiYyAO0n1fjymWtPCW6U+9QS3XAF5q
HZkv11VYyKA2rT5uPlPgiHfZw3hF5JVV4q2cgFRMdY5+T8qAs9MGWQILfQoiRsdkx9CMuCHRUlDt
47BVom35liAXhvNf9Qbamr6u6PIvpmHCPjwvHHbSWL1iJvo/CV0tPnIfaK5f2o7BIIm7QOqd+fSD
z3xet+EMQ08ELZwgPXqkADT9mC00qypk9kY43Fw2s+vDOdxb4pvvgWIrfSLr2gpCZCS30MEAP1ZZ
IiFHeDZ+7S64YQWF0/XapIFzaMN5ZwxuZiDm/SEZFkUaCWuiSc+FxCpnnjM5jZyrJqY3zb+UJ/fk
zjF4u66K+xv4a7UivU3q0TMIJfzAd3MYcvY0yzDACJr80JMqspnGmvydK9gM1dtfFia1Eln1PaYf
kxOXk7O6bV2FoNvN2rXUa5sRxQhXE0Z/RbkjN2pk7T0H9W6juOpIeZ2P9jyxBWjywHvJHwks9LrB
djNqd7VcCmtBkcZAZyw7FSUl4XhuXqqevblQew21fULvHyj/4R5LPmRwjhulGIqG3GenvhWjBLJM
BWIg/tYVVfcfvSmksGVssEvoAJq2nZgpWLTmacg9T48mkADi6sn9grvcYGkqIBu6QzWPdQSgs2/K
vQenjEA1T3wENYZJdz3tRoXeEynCGLoePRrk7+KSkWWpYjRKdB/mo2PTaSiFJq/5lolQlGV3UAbj
RMgFIS8iC65yRVDr3FeOObTgvoKXt393poeWob5w8Ece0z3Wk5f4ia3lR8cLRf4zIrDxJH4kRU7t
kPYeHKD0WGVs4Z9zqIDVML5aIbNxPzk99pgj+nxgnvzgMZjHJoG5CQMZcCsDZ4T2XvN0FOIzuyjY
Xc6h3LmDVGtkvgi0YAEFsdJFYOQjktnI061ZnSNlPe4t0GLRKyZEnLLR6W7fJSc5yC1PT1avoUe/
dccWWZwm2v1G+4TTRQdcRne7UcEFL2ocgXr+Jy+8azs9vN9tvQ1tBJfn3R4gCJTPOwAAs9E6+0qd
SJsYaHQs/4gY1tnikXK6hAS71F+oBt1HdYpmqrzjFbbW7O7J15AfqVOHDGN+ULt6gZzFgvQGyVUu
JmEf13HeEMKyQkfd85/Q9UQTOWbUxwII0d0ePjavKsIshODKaj9Z8eqkSWgQ/CQzZ4GHksEcTTUS
4lo7nKZcB4z1TVLNA6u0EDSmelL8j0M5VcOwaJHnaGGIEriOEPVHnfHl+pEQJtVLatscXvT1TVF/
h5TyT2T8ahSuvQiU/gfXTyBKkC2d6MnS4MVf0QdCsIvG7sR9knPRbbqSoiUu8NsVJsBbgVdK5qJK
I7nVLUGQ83FsHE+d2UQB/OGQPvJD1DtCORFh1S2Lk0fYV/IOgEOMoQQ8woU6k50380Jkx+XaJ7wY
4ihGHYS8Pc7OdLEVjtNBRkTrb7vSu+yRNBHyCt6E3A3BS8pgAb0Y+MsFJGA3WUA8ZH9X8sgGL0+4
JKFDMKrIKQAfNAsTwu8Ay2bfcpgiVAc0dXWoSntQuTIeL38pXhmrgr5+LmTOPhIwW7GW4MXZDalF
L/X6+JUYPXNDb+O6ZDPaut42iw16Caq4nFSgWKJ5anX0j0zjgb/TTbCIBP5gh236iza3EPPhVe6Z
Mvz/yu9AayleiXOU/KSgK7Iop1AOqBC4tBd06oDDodAbKdv65nXiVbwp+h28i+E3W9ZGVglvW1ZR
lnQf8fuQBvKQaIpBL8EHGzFdR1Gu0KqwNRddm34vfVe6ih4tTYqXn9uM+r78oprPoB3mCmFjQRn9
gsVqMlW4P1LXjAuLkPIlwCm1Op+H/mlxANpDtGlg/u24sHAf7qL2ueaEKiJvOs5Aekh53j3Zynbz
+Rq3TmLokImlhpHBYIKCOlC1ddRRcX8i20HIlg/EE4nunAHVFGpd4ghj1N8XfleX+a/QapkqSIiw
WcBdY8nqbVcmCXxrJorbWoCKXxTgx0KTC8hDyYQReVsFRezDO/8gw/9qEPdAqTbr37uN7yIr8wL1
0yX6U5ftuFvWSZFv8q0wW97TRVu4pP2y9DpcA4In+QrDw882b5n6kdoF+1HTK7UahEQgQapOQpTx
ELbLV0467yOxHhf/V43Ulw/lm0LwWcXkjBlZeM3CuYfJpMZgHlUcVM3znz7jvwfE5QYAl4PDxFpc
0pWYpgD2Jn9I6U8NmS7lWb34vIjNn4BfyMTGhNODXkxiBRddF86+uvZJPFTQeBpTag8T7wI12YY9
r2Lg3LrwTPN0Ja+H+S0ETGO2TSsoWQlhRgJlofGB3LD7G0g/avGCdX+vvbGaIbWAuT2ywPhTfNGI
KM048Nc9YnggCX3658vPq2r086Xf7DvdJwlWC+0yZOCZyvprjoWe3rPdZVDoijTpr0+yHGbvwufQ
MywJYnxVCzHe71R1dTWTaOxuwZkmmqn6XuqfRxrkZA4LqhG/Vt8LacG6Qnu6et7u7jlyhMbV45Jb
QLPUS3/TgZ2xkWhmHMrRG8j40dD7R31guuDVhp3t5Z4sb6+7FCUJAfaHyECKu9wNlmr/ZsyOuRh+
N4RL/2duZXkSn1BbIdBiUwpM6mOQf6Pnvtndt+ev9kk/puIBAMZHRCj/FWI+euIqTrfdSqRoC8JZ
ClYV3XFh2ZlnpMk42KzYk8ULn88+ZNE+P8Q4ZpSXGYEbD1v0X/A5OFu9RaO8xTvlZVtzGxtI6kQj
lcYx2s1NB0neicldvVy0CUvNpif5e7IsL5+DyO1hxCk3yn8Pk27I0uK6b0mHXVni0NZz+aYWaE0D
T2NGQ97hXz3T5vbugISKnPbQaV3GDlx4VeG2/o+7Lceig+yPQy2+ec50GXZk37OXjvavdsHeGfCF
9j96nRGEdR47q0cY/npBdFh3Fwdik1QoqkG/+uCSnUfOq+QI0fC03XJDcCJWQDw4TVmy3tA4j3us
DOoJMNnUwelBiBdodma4GSitj1r8hHFi+nsJbiq1/8rvmGPlLdBNRHHwtf3IrXCk6TXRG77PTav4
A9VSKhpPg/NpF8q5719QCQqeZ5kWjPofYX8ptzYHdzZWS2cQciOrDObNaJv+TRSD6HoOoRjzqlzl
iWekI9LKtWWiErwPLqZjNnJ+WchOBysFJxc6+eK5JY9PZfnrTYmO2S4HBU13AGrGna/L05JKPvqt
Uy/YypX8b4+RKrPW0xgeY/gWCiABz6J+MDnWL1r7G91EPe30ksL4VQLvB6Rz/3lKTiMO9qom4z1Y
fQbKoWWi0cxHLBp6Mk0T15znGaOswDPkMJFyUR+ovlQM/O1WVe4Q/iycOkCP6Tlx9jP+zTemg2cj
ouuablUuuPPn19tBEJpdlRFXD6Ah9p6VHgc3SjT6IuwGAhUHcGBBFWkPFKWAcmxV8Df5op7HEhAG
q2vvQmf1IXJKfjCq7C7+Qsp7FrB8LFFPpUmzoCy7lAS8QCGZ2cScJlJ7W0fYaeOcF8P8GJLrFZAV
zSAQ1ynu8gVXedPuPxqzs0esNJ3x4hRxqfykupX4PLhLWp/wUOmJ+a/Yomj6/xNZuclFa2t90Ime
o+xT3RiTdbtks091N/jlVhxnKrHw63jjoKJ7EyiXo9OIqMja0uc+7DA691IFodWqf0n+o0babuPv
XCwyD1/x/kZUnTCsBJOD4Q8WqayccxpclmndanIjOqZP5WaxrD1RPP/yGY7nplplkCg4Y5Pnpekw
7wVrAXf0piPN7PfhgyCt/9E95hLDopLaSG66GgmkkzuII+e9d4R5KGricAthLoX0ZnRut2EMtgq8
2GFixb5yMlTpw4FQDUi60BI6ZYFuSZYlWY2cyKRefa4Kg6kpd7v3iORg/DzxnISDr9tHv60ZSLVt
GjPGsOT2AVvG4rU3TFrgcjQeliMiJ5NJjPTFDFCTASy66X2PfdbpATm7/o3SwIPYKtbS9r/hNoyt
rGguH4xDwQl6hGQMU9kHMcHts4J5D+OtInv19DIcFN1jIQuVW5JfWSTxiuIJEQJgATFTAeAkyQVy
8rGnU7HOC4JKdLDpHR4c3APQr4k+93WkA7xDBuF4eO6j2jcrNkcGEXdt6VhYdkPcS8omlvw/jLdX
oWBXcnaiiwRLLwn3ouEuBtLpNvhiKVeelb7yd7+YLDyewFggONIfZJXnV+Q6Gc/hhPs5hjDFSztl
aycnHE01iM1UgYmU2o7Wiay8NTQHkKfPXGVmtVeQ26yW4tovRl6JVET0dmRooFoZd2xMorxr6afp
pZiHYB7RWkF8TUjMOgZKAR/8GMxz/kPyeLriO71bfRLJLVaV8wt7dsDnAo3SRkffV5Ducp/LarRp
ZF8XvhWzpXHDjsmHyhotqFHI3r51Z5AcUwstb/rFXgC/oFbm6+t0Nh7O6FZdHElotUA79WO9j9sV
I8hTVKlu/+MpwsHBOMNJx9sAd/muyf0YqpC1BPRGPowIdPtoIvLSav6/TVFcUu3al/MaezdbdYF2
kudszG8bvUdEW1GiSBEOt855F8gdYiaPGlRQYs6l8vdgdwyN3N7tZ15uoqoKgSKIHy1NfYh75o6r
fM9QEHM2vi9BnG8BD1dcyLVPvtCLfayE4BMDJ6KveZ/Da9gksoJX6pFHmwNmkrPLaYdZ/ZpuisIP
g0JqaO61YOKwoDmSRb5R5Clmn0GksHyBwNQZQfojpbJRqjzwdT87DYXVU4JL+4awinEUZoHkvMVf
hBU+OB4VB1YTsWkSq46qulA6FBV14O6J88JjaiCKlOJ8AwGtnNs/yBgFkiGr9JoZiEPWvfBA+TXG
c4AfSgmM4hKhqktB83Szw3ZlaEg6DXYqOUWdEeygKv6p72JLpVSZ0NA2Bl1pFuvnIDXBAJlOA7Cm
2z9kNGG4GRqjZr1j6itfav7zBiFpdg6yOzpyw1UxFgRxS8b7JkxyQQt+f3btSbVSdmja0dXx+rzq
EPadcwxQdwsUOHVS28AFiJ7UKyKM1c+ymPzO2GWL1PNWWjVcljs2MJvne4MFt0/PwvRuIfZkByic
QwX8+6TEJDXSEfeRf8icfmpHPtFC0ohdCfJ23QkCPk2RBgUwXd4U/dA88A5NjshxdU2wXRVYzhVK
XU+Cx2E9huoDRnrjanJ8Wco1EJQY4ZIHJb0922hlT/ychpxEM8DA/fZ1os46fZhXzOG77+i9bvP3
Qe/pnP6JWv/z36EnCk8jekO+Z271X309IDUkHlxYpePHxr1FVvlwJ2iHJCSvRmUNxc3nw1PVbERC
fYwcZ4JUs7Mu4axRIbSPwt9v3VNLeUpGaIlm0woEkPd2xj17T2GlS2+Aia6jcsOR9l2WmwkzyL/r
B1DxawqgXU/yrhYwykTIuI43llyWruJMfumJWJ0KbZX7ubaur0nIDIY11z9QAt+r3tlL6faFRTip
A6GLb+lxE9AJNFu9pEzWV9zIhEhdCUNrQud5F5i97aLmKalmbs8MkNduOR/Z29D+P0JTRAh5fNvZ
J4y3VqyWNj/7bZgVOvrBP9uMB/JIawXoEYBbLWv9b3Ve9KPv4iB+LvCLKt7kUHZzpnXtw0WbIAl1
01n0JnVxq26VLnWzm/xbpg/Nf9d/Gz8z6g1rg1QzzALBh2aEM/FRrVPurnzJCgG8Udj+x8pXgDvP
UDjc//MZM76jTds16kfeToxKNj1TcyADRE6SCIJJ8JTnN3AGAuGwoo3sALKQFkAKdVcltdnibzEZ
CwuXDmBi5wDDvT1l0PQPcJ4n/5cZxwJS181WfVem9oh/jRWgVzH9E1XJNgTOEyLfgjzI2P4QrSg1
WrVgur6T41CIfzYeet+BgFsxTz+JspHjjxzuEqIAURrMK8LAs8xo0B1rk02A/A3rGTXT8HJB6vAj
IQjVlOP/Ok5n1Ewimg1ilQuWddxjEqlxNdEFRQ5ex+lweZobuit4/V7NbZKPYn3pgDVSPqO+RGF4
lUj8XIgyDqI7wh7rDWFYhaQ7e/TJDEb1B4Zzz0r/EDLXkdQrP29qLzeot1xGnWzT6/2vOyxKhawi
3amTS3XzeqAwy1jVpSNrUs4hmJd+HhNLwQp3qeKHiM5N59Dod09T3vtMaApzf6lMACaNZgMTok62
6ySqBrwskFGa3oUtI/rMHNQkOy3ma36O/GeGl1/6xpITbY6rZFjoIyo4ADHOWwW8wU8Sy1OGt6tQ
t7+VTWAlvD+Yl1ByoZGO6YZhdLMUhzcjwdzJ1h4PgYTPwx5i0tDHpDG1bLnivEZz0e7ucuR3YM9w
ZrR0LnXUxZBMcdgmprrntzuZ/kYD7v0fWAjPg4OJtNs3RWvvIF9xofKCZOV+sx3u4OO5ycZIg/8c
jCGMEAlSA9b1tVm53gogKUfpwTqoe/2sIQr31j4eexqGh0+V3iUkMw/E2WtOWRc/UlMKz7EmHXT5
6LVnvuNV+8f/Q2PjqFpY2UCz5dYaGHZcD0c99EkPuwy00a76mpjcsWZ8xt6adN+TXTXUjvyoTWcG
PHZSn0oVO7KcrZaSh3if0Br6LvbPFXsUjWLLbilKoupZe+rwOVnV52S4LRu+kbHdJhJOlgzCGxhf
FA/lqtErgRtq2fSLzwtj0tivUOC149b5rBHXs7Te1p10JqtSyrJeTl9QzVMdfxO9o4kLacRv/99m
ZmvTtTciDpKl/r8Fb6czl6Yh//lJzboiL4DmUJsE2bT9mBfydyTfws3JZ2WKu0HvFj0ceIiCbhdx
h+Qh5rXulCCWdFeELcRujfPWM9krN7/3eHYvg/wFfRWy5tI58prmTo/fVZ+HL9juQmF7Xhh3Wrac
7tMiRx0nH2r2ZYKktVr65/JxMXVnSLTYB+2gAGC13CvKWmEDNv171RHLyHxw33PpPNcnPq0I46tE
akmCTHsacWyuDBRW6B3IKpaEHEYakFaBIn/pJ5gGqU4ycV15h1hmfP3O38kRlVEqC001wApasc7G
GNra10E+kvL6ms1+e8NRRxUwFeOly8aILGHoRUI3LOzGBsV5eaLVBND3JaJ3b35p8D+dPPhauTcQ
EvJIGKCY3VsyEdof/Eyg1/MlYYa0pUsRNEpB/P/V3vagSt/VMPfWYvTym3nRnZvK0jn5QUhCuJIB
I8RXzhA63hkMSvdrPmioef1/9BmTPa0Rwxuzvym6xKl9YfbSTFozmLaO5izaQnIaoj7XNn74PIiC
eJel2EJQ0M39hblCOs/4S64jwG14rwtUcYrZtjZgjKb6s7VnXJF1Tu1/C1lgTgyZxRKeLDYBWBu6
hw9iHbX77f8b2hu3Igi7RH5AQZAsIKymV7jAqbcMvhbj5HvKFfvBX1vWQLs0laLgLD6ExG9wwaI1
dc79muv+coCTinL7zSOQaOyCy0xUMR8HG1JhZ7qUk8pP0g22t3gkHhAqwqO3XBXym6J5uVHFBsb5
S+/Z/tvavH/eqKd6gVQdF8Hi4o58y0U0aYluB1XiOYC0klgdEfZ2EeQ9hyRKoE8Rvh7O0uC6gMlA
c4EUH3YSWP+AV7esmcxlVrGdgWTZs4ROZRgUn6XJ/zPvcvUxpy9NcouLKXY34umqvhIhcwjQ/aaL
bBHrV7Bsaxr4dSgvM1ZxcvLZAq4aCbYE2k/zAEQRrjdv5PqqyenjdFuewi5yGQh1s9VKtdcMxo2w
6AlJMXOB3JOOCBVInbSYvjXv7AKGHkjKWYTGCf3Mjt05xfI8KwUpqF+DZxFYAaTintE8Fg7Rg00n
p1XO2eaUhs4ExIxC/z6r2tOQQ0YowqXxrYO9JIZXebdPe4XJNwl4KqaNgWWDH4URCwMY6Wxc0YFs
r6+V932VVBTAclLRXItuiDQGTiBo4QP4+uD1KSbXslrQbr28UIJUqzxIrBRXM+x4O+B96ink7UFL
IuV95XwsiOwdDPiCP5EiD83QaUkvMPsydPeQTTAW5ONjQL6mB2qlqTJlo7RrH7vrj5/Am6eNtA1F
QbIZ1rpkUvTYr5wVfCoDnVmHaK0Hg17F8jztOTFZjwEz0ncCOFNEz9qx+zyb+wp9offteUFcP+eN
DZq9nOs62VIpdulJ4guc2p6583tzAyZhSBvo1XiuiJejE/AHOoTHiguUdtClE0rsp764Zl1aJTs0
Lqdy/ZYMrz05UhN088BE6lcCkWDG/hAP1XsQzR/CBS18DkHeu/rLmsiP5r+ubKdNxKJzxE3WLl40
j6Lov9e98FWT5qfJ6kpDkUPnN2AJfr7jQQO2s4hdhEhwI631s18qL8kq8QOQEYyykOcGp15j88QI
+NHphtBCDnXTDuG26hQufHtQWJ4VTLeniXw0KX5m/F91viKUl1Vfn2BtFBn2QATEad3nFHaCBLx5
0pEJnr25bnbI8p+JPZXYSORq1CExgfne/bNyHU+wOkG6FCz18ntZ+6EFsrh9nS7k0B3iYRXjR70w
0qMBGqG1d/8ATWofc29dZIXqE9k/RZ3IlicBD6o+8dkXmlYpz4fiDIuH3Uch8UAR3PrQXsAfd7zQ
psZ0U2j7gsc6Pqd8uJlXm8rKUTp9MjiXjmFev0yz2TPUtBG5+0ThvIhwVCC3ySQuV+A8Xpq8WpeP
3EKxbmhoHjr0PoJmX1rzheHkYOIruBtDCMY2I+/omKqtx28VVzKpSXNv0qcTBaGhPAytS2h7VboS
wZGwZFq/h+XxlNqW6V5AqQXir5GfTwhEb0HR4jrcYW2pRWm03WMvK+o9GrWuZ2bqmIc0eNP9D/aV
mae6r4RQ6ZNMzBzDpx/8zAF95gt//M+OWXYmm7/TTsw3lxZh23Dj2rHRQwcF4slCkmdDekpooSL2
QcXU01bKou77TC2YIgAHJIRv9AWdciDTxJejNjpQzq/5S9H+Rn1XdJdyorAjT4I4vF6qdY3PDD4p
ZbmBx8YSdc3r0wQLNigls9cC67BJtToxOu3Ft0AwvB+R5fLPgEmyxVqbx/ESbLaL/oiyFJzxTHVu
xWiMVunD+/wKRbEasdS+RM4zL0RQzZ62XyHhsCrAYnYSnRhDMOwMijAW/2RipDzam3CxZq28oR2c
0RuEarugR6BxRXoJo4++R5d6Nt+TDFUuvCKC4MZL7j76ND2v8Ydd56aOI+ei5B7iF34wZ1ChB7j1
vfx88HgIgAGxJz8GSmXohZAwH802V29bYepuCygDptHVVGVyIaUmusr8ZxputeiSSrsaILwztY/u
fOCiY10xLhuYnqCzNfFiXw+diSUIMmv5YneDRgp3gxfRSyvaoiot44DtGw7d/u3MlutFdEB+Dr1F
ddmX9UcmK5EGK198oWXMMkhlvnPpKGiDXMwDPErxE/N9QWsgi8M7kvoiwdvFv2TQGawAXeEh8gNn
gALO6gL9hQMWGq01ga1iMfO65vpv1wjibcuOuJQexCTIkmzU0IRtXmtKu/xGVICA88jpP4FXxWRe
mo1w//6pW98FetQ77yPht3fDz24aGaTkQZcnZkjT0tLX4tVCAgsIsXjWa5/Ono7PBeptWa2fTeKY
U6FjeSCSOfoljzl08WNDY0yfEClbVuljcfKT/4aI+PytQfVki1gAf5OrW4v+ykcNEmWmRAV8pNDB
aP8gB6DeTL6g11FhGGvHoNPZxlyejeepIInUCItMtAXjWJQwkf5g4B/ngV5P59G09vgTXWD2H/ob
GYLMZI/XYwivQsQQhJwM5gYPTy0hflyrszV7A2CtVdeYj8YsTBAgHtotUuH5hW5qa4lwhIWrg9yX
jlC2KD1U9yiYvAOE85eK6EoBpjUhJJOaUXaW7wn50vRQXmna1E+MP3Mk44UseKh0YmYRS9T/IlA4
0nfjNXkX8RU8y23jGqIhyQ4qSW5utmkTnCQDp+XvFenzFlKjBYFr6z5SZg3E2AsFjzQHQJOWUIii
iyax3aKYZ9YL7kFY4ADyoNqWVP04ZajAsDsNff4vwiNNf8h8lfNFivFBqyI88grDFbguXZBEojwU
pv+hR4DXSOeqm1kqfQSL9cgHzeWbONTs7LXWJ2bjlbIsAZMFTRFT7OYx0CVmeNX97AliHzlm6EwX
Tdx9hjpHtlOd87z+zfDAeHwDMzr+anTcq+SuaICsrXsezECXAWM07Nk7ysHhoF1Sdth3nSlER1Qi
TQsPG2wU0E1G+Z2UjzQsZ3fMwEkJ01FFq1l8kX2XTry+1Vok42ZQR1QC0uvzQCnZkR4FczutamL2
DzJAdipMobYQq92Ecbg4dVsT1tQsKE/DI0pEHIIDOt5vstkvRxR4LNwnhYZL5kTC37PNerCnnPaJ
IjKPxcclrAOxxqmicrSXq85NlzLQe+nnECd4j73H90v7L3NGV9Tj45ZPW2ph0AwsoyhwtNCSP2S/
KNd7Zx0yiUKZ+sgpUgr/lQzBG5ECUaI9TugIR2b/p/+6u5aLyqQphparXswHhPyA41FUFeAtQPVq
c5gDfdES08TFi9v39vHB0daR+vgIdFz7FdNk8rUuUDyVKYzGFvSP+7Cl/EIlZGrurmzmg4M8EdOI
iRcsqpDy3uKiI2TosGB7GFwrznkJEYmhxktZpEdOvyaS1tRd36XYcLF+ho60yus3Ps+V4NAT5Qqx
GIRAw7rRlqzEgLna2K85GKqgxGj3go1sax/qWDuRN5ceG4y759/zcQNr58qYrx4/iqeja6vuh1rF
S+ns2gSxpD71w1vdJQQGMf8jwRg7Ht7pxtNPWjHzxvwTXoeegJKtIyKKbxpRiDrc6y38BWb3ZvoK
6wJoFpm77KuvhFRkHFrUvB0yPh/ORO7NrShvRsksx9iCoDh7RIoHQfJDojDo+MSdjfa72982esh8
3mVV0JWWsoRYjIV5AYEMdmIt/wnaiVFoGvuRq2OKL/eU662+677ShIQg1yrZWfdY/kPywTMNcQcQ
fjcbMvMnSZ4BN0XTA5aOpEGuelcLjYu0/ThLjP+gRz3jY+4ePIwH61cvYBomxYOiqbM+XUvObaI5
zO76gkdJ+qWcLQnUvcbdkhWoSw3N7n5NOiDxOJrZOvE6gtit3BAosNTXVEKZpySFwr/wKAT9jlfB
darcnF6JQReU94WRW1hsCNpKXZX4NkkEeCd1Ggf+rD9dsJrrnqjqQQoL6MFqF0FFf32N376BBnYC
sybSB5H4CLfeN9a4Ty3Tgq4rx0+tGBjz+w2apuZsAyXIY4z8KtixRo7lYvh0yemnUlrrJm2qf8xu
RmWOlQanjRQnhKXy/M+wNzEvlLs/vFQCpQW3uI8PXG2JlPWh0QjqxJPmybwfWjEJ3Tw+0tyQ+SZt
Ql8cNZBsFC8nRZH1IHjXFPD3UVwZpX4gKrc22vGoYfcXxmlLjWKuKdiN4M41aQY45BmTnorRfTwJ
WD+HDNUqYyJDalvh+B+lfNUM9krPTHJSuuGLvOZKahV7q6OybwdzSppxJbp5sOJi53V7VFpYv7BG
Sa5OzYOrr9JC1jC4qcAz/uMBMPhHq9PfXI1tdzRgCI6RL5AGeSXhILQSVuWdJdfQfogmsNQi19/S
ytrETVePSL9foCAEv3Jkwl7/JE7omkDydANjPpfmoKuFNATbTw13x3bCrkZ+tSGQ1lcMUF25GNGd
h78mw6bJwkh04tmlrfRc2Moqz1wav6ZmxsFetch506mA01PODCBtP2+KYtffAHreLGng05Ck8ORr
8LDWQ6f67jZadDq7ev/uPr4zYxZO0HORETAuDIVB2Eyc3JeA+htRLnXEAClxXvo4kdiuvgLDk1eY
xyFp3OpuuwV9rPgH4KcbDulPw41oQSSkNYMraA6MGf6qYW+MYgp0pZF2MSUsv7rn6R1aIjpCQCCl
1lWBBVVK8zh/004n6WCDmJDpLN59PyM4XNDZUZBIG2ebz9IF/ChVbxLTKg/7SMRWXHNTEHaxyXaX
3NXGOwLFt9lPi6Sy5P2lEm+U9o1Tle1XBPoxjm7k/JSkoceg8F/Np+RtpkgfqG0R9kEQaIvyv65j
bD/APK7vR7Ta70tS4QTlhQZ+AWvHbtlhx4Tqkb3GS8pmRnxVEeo7ueYtRSm2RHkFQSltcWaQIORw
QHjDEaKJzLyA1npUunXDHvwMsYQvEI44M8/bj8eFUuf+j6X7tqOOxDhHwyQC+T4QvNwYb599GezX
tRZMTGc8WJXEClWEmD0s7ybgEICtKXwpPu7EWFIu6k/zs8/KqXTS4fq9WfyUCK68vkvONB5A1qij
x28HydifGn9qvV6GplCm6Qrqrug5GBHjvZVMDSxxmpa5AvliRKoEAEDigR3pHmasw6A4kGCocoEV
7zKUxcoLpuzZqSRpTxbVk6+dcLbU4IjLHlOcDfWh5JCFmMSJtDXKcv8XR5Wk8DA/n5PctDG8YHRP
z9LSiVH2pyU8XO+ScvolMIHgqsV5bl5scW8kPpiMrRBULLcBli43qL2MWqKIUFm63hTBMMHk8Yp1
8/aRubxqDPUnPpxqQMv1nqe9mHgC26aHdR9DB/PAcECueudTACgKs0Es/1a0lW4A9apVqEpplRPk
mAM/nBEKB8e4JQfDZ9BzJVQeKh+OZ5evCHnHS/tJMVsWgiUafl3xM0uHz1e+mGP98DKFMQtG0VQO
XboDQvqRPlasOtL0EAVhA3qFXCy2bZjtUSp5BDIK4nq5hgVkrT1rXA1QP+SSk3NLnb1ltmxZo7RA
d30wMTsSYOpoD79EGG+MUq7HwltcbpEQ+4Eob+Rm3yPBtYW96fxp+l5pzr7Bf12e3dbwq/RTRuKv
XCD3oy/9tLtbmBMbuqcz8ZA0qEjh51OGLRQnyQ7VYBOghapl+hvCUcbgTTAxu6AwXo2m4x3snJ43
IVeXzRnzwGg1haZxf81hil5KUkc0fpquyht/jtIoS+YSyBsVkrazVDj1naPKedT3VA1hlvIj7PKg
3HVPM6rwUv4CcupT7dhYPCl1K7iW0SZ2Lb+EdAa6gEPoIGp+EOa2NzI9Ij53ZXAaOaZMb58uNUVL
ryVkfO6RgEeTAHAlddGmlPXmqa0jzkAF5d4YwFPByVA9w+VHZn9dVUXxSaPAwWzKp+XjjiDdOO/z
VD1kFuqIMjQod8xcoZgYgC1Rf9/uIgbFSAjSHoewwCiZpXkXp0xmMAkUPsofx0l8GpN3kJZl/aXh
JWrrLeusyZky8iCKl6aqA44lmJ0TMXMLVw4C7kfbpS2dc9t3gbHxiXCOWjuVPDlNlfFzwWDT0/7z
NdHXuthHCzmq4rW4p4OKpuLjAiCtPPhYng9JgtfrRDa7CF+Md945qkDB36ie3BTaa/CW5PJgHYiC
qDPph8AEUtccxyMMDA8Q0uPx8LrwVKkaqVV4gKySlXXL8aW7mMJqmU8Za3ucuaX519KO9ihNfgHC
n8OJD81hblFJaDRlquYr2CpQrM5ba0HVBLWgq/mhufofw19OGXyHPl8NOcREcQsFSCzYLrsVUojf
bSjFCfAquu4Y5XDHgPDuUZl7tpCcUAORHZUdC/Hdbn6GqfxjuFXtooMywbz8H4lKTw6HOK+6Prp/
45y+jjfFLK1YfgAcPUiPFb9JVdUKgtBIoEm0RjegJIhA7g6OJKa1fN0WVTSAwCEN/cFUH7yeP5/b
fKcXL6lxO5V5gFHfPzx9xkvdBG1PmJGWQRQvVwDIevO87eVuAs3bAfmGbf25fFfWuB13i4TKZ0En
/aXs0qJREegII226M2+STehDIJKvphipjNb7dz6YN9SWUTc1R7iJxSCwn5OuCiERcU+55irZ1tHP
fhcOgewNqltkpIXc6YFJBqoUVb7B24e96ewNx4vQDC+Y1nxUT7GpSu9KKtxu6oHV3y1xvhYHggfa
KuItmXgO5bCDEqWkdgx9QTJ1hxAxy8JuTWfR7PlOfZi5SiTt32N0KWbXvX/tu9U6PkIqkdtlmM78
9fFvFg8YarZN8jpLQfuEoTcRk0/r+SJZ8fD8tK2+M2NCS8HYJEudf45F5H7YDgWbPKTJX/Qyh9z8
gmwoSnj9uq4V+YtU+rDQPGyvrJRhc8iXm7jBdoDB1Ct3fv2UjMycESkVtjWX11pity/wntoFGZTQ
3doqE5koYD+uEqnuSRsWuuA81vZ5cRYbMnjM1ohoQJ9jCrWPIH7JHxPE/B1Yuq8jQh7fg/aTQpcJ
dUjztfnxDj4tpI0tcyK7qcaLzLfYs0xEjMNPX116Xjq+YFxdbjzhtu5Welt2KIx8Sbzfh2I8qr2f
IUozG6RJvLuYOmTN0Jsb1g9j5Of6THfI93srFVRoLaejiGQcuuRQWOdF1Bpu2gmADOkGx9dyRkYb
uEeV3XEUQkXyspnfNRmNIyt0zu5/EJ4955wR4dO7sY4ou90zDWa/FCyy5eNSs/y3d6xAXTYrjKDY
WXafKvwyQ02okzFXjDmgvAkA0Z563tOBPyhhEP0CL8y/a3tMqdwu9TTpEUso4Jotk8F4ZdI+KXYi
dIisunIIncdnhL13dl0GIEnysl8u5cbV/uUdCd22lsEWsfQwxsG/JJ5f2BJF5WfTovpIwdBiHuzn
/pRMsIYsx+1W07BT/7mbi5XApBZQ0EFimDEsFlxjQY1IQxzVtCCSyYSJVYPipaikLxJAV7A6oSNZ
o8DEl89xMxcDHsVvb2APD6TfpegSBKtAA9zlLLl2XQHZ40t9ZOuOEFWJHUwfz3ge6q6DA8izfYQ4
DoIeiBAPcRirhw3EAWGbfWnGJMkZIb2oUbg2v3Yv9ZsbR6CfMbItaJP7QyuR7XiHbFxeUqMfLDaq
KQkYmc/MHaqYPL9KbdpUZ6Izigdpr2M+o3XFlcC7tsZ/nto1leJgMR86iakvFgXojvONV5i5F8nU
baBGHCpSf7G1eoP3+4YxQ1l3WxmHLkrNHtDmVMjRYry5FD5J0D5fA0jfyubo4hYY4Rb6hW5Qez+o
35wPiE/HDiB9o+YbfJqheYNb+eKrxdWNOwwcgobtNlPuljgWghijXFzvSmhn38cjwMo8vmoEqq8E
AYkMBAnY5VQaYGXvpkz26QX3uJyePbaR4G3SLtpgItc0+XhlQtnjn98iYzxq+84wlpr4r2q9hXgJ
/XYNyFkqFOVDLYMk3AxNV8y1wdfxDHMNx6gXor7O1LWN3ntzbiDYXudayhLX1VlX0kxXOjj1cYYr
OStb2bqTwPjS195dgSib7nJc0gk/W8wucyQ/Duac+ZSwn5/PRGMpotZKF0lPLrFOfZmOey8S7kS5
Hyil8lBQMYL+OfiS8CNhcLmtNr9BoQD6iikBpxBZ1sR/WM9dD6bvtLRUwNwEtmbWWZeO7iiSy3bR
onkExILD6h3WIn+oeNMzQ7FBNE0UvKQQdKOYoBrwXwx7JycMFF8Ye25KVmjHJQpblfCaaZDIcAjk
pi79J9ZIYRxsyWRWHHM7aMFRFk60CM5q7c5jzLW3j2kV4eevwvSP1hWCJ6TLdI6PlRubnuhGTBjW
IWZH8wObapTaTUqOo8WxLH9ixkPzUxQS5JjgyNeU6Xc0wnXWZSR73RAZVC9KtD1oJJ7TbAoAmPxH
Cs2v/SFQHBQSprC03TtLC6tEeGhMN4Sw6+15g9tx1vt+KXU9iqvJMvLvADZp4tdFJawl4k7tu2PB
b4D8r+VTSNISeXwkweAAXZPdCxd5Psp5A0JE7QufpesZlzMbyrFYoKUzJsGXTW1Jo3IE3mfY4r9o
+O4gqRNulrL2ZM5UmwKv/OffQRC/yTFTKWSrwBzxJqqxm2Q3FzaKR84vl8bCIhPdhWwYqSbXUTaA
mKgljtgHaxO5kSksovt+ABUZDXFj/Z369AJA7IjslaTECEb/H3wPEPvTeSCS2PxDqKYgK+slShyB
P5od6BCqjFAmEt9bZJakD8TQ/Be76wh41Ht2d9U8fUNQeF7tCbwyrVSe/lz4oLpjWRJYi+RKW8Sq
scRasLJXX0fLfYZQXi0VPIJWGJ1Wt4Rn0S4/0tGQjLx/rCIBVkNWUsD1ZcAa6SGp1UXDr6OLNUDv
5F5v8ZiLsDwvoLHz4nl9yGb83qmWXUoe57gBSDDjSWoBUrCBb1gntwoy/nNrRUaz5/XaiPL2FgF3
FCuJvQCQxOjmNFWescl6lK/l/uXHlK01CADAf9fBnpNoVCDbxG+22sqBWZrS8SXfws1ZpuqWoP8l
+3CvYzRfGO8S8qRKExObPcN/oMATLtjkD6U318IIYpVmSVqTJSwD3xejBOPXFf85q5UWPNK8F0Qv
zKjPoCcbIL4pmjyCFfF778ii7qzvn86eapfvfVFrIaL4wCpti34hXz3JNPODMJCm7Qvh/lJ3nFJo
rF+Qiuxpx//PxHwUr9sAPFaW20OPxXTgCQG7uusLQDhSwr5kx9lq5sGEQh2g0M+t+wxJU2wWeL2m
Po6SEumYUCqM9XvEutKFxkZEfX8URk8iEkL941DAPjKbIQDcyB420ytvnoVwLbB2viMGYEKgFdEK
dOkKqeKv+eOBM6Kt3xmeVzWBijdlfYODW58rq87VcGiL2UQJRQ8EqYxBCvJAsKnadTIuLCZji2HL
kY6A0bisdnbbSkxJ8prhvh1HDtM2NvWO3D/gLf0q/QTsbnv8JD2Pst82T4rkfLcxS1A9THpFDO6d
iYMLzSRte8VI525dnmK6yJVlmW2MR3+d0rCxctHp5rqxJgZWaOv7hkRe3vy3J4+nhr37m0sUXyOX
GrXnhjToptwWu7GeCElkV8gPmOWHXHAqFIg4zLEaxizs1kM5hH7yXgYLnSwTh3jYrzYyV+b9foX/
cAkEh91GgBQ3o+XftKQ58b9MqupOh+e70ukoEmsWhzdEbyKBsfDIr6ev5bUKlahpH2cuiv2ltCbu
IMxMEZ0imHkxPdoy4+V/AyfhY0H9FgxFns7YA+Pz0ez9GZCIMQBsIsB1Hh2Zc3kp6kH7YDPT441u
T3kYdFJ6WB31qXPoBwjaD080rPnGpVy6+GCo/ZGMHVwIqUc4VmcHpaLG636DBwCMqGICRdlfbZp2
yMpD9H2v+xCB0M0rUw9TyKgPAvn3C0HCKUEdLpKvQBw/WRQ+CAcIoCKkaoV4daNUzcz1VeGEXZSQ
iHxyqde8AbJassAWH35do4GecZY/gbXHvS2XC1AzzhR8t2eVsfEDlhgJOM/m9FmBO3FpOjlqWNEl
6LLVIs+sACvNYuHOcJKD2jFcnmmsrVXerNBqIlcb4lyLG1i9C3CYzHO3TiU0N4YoxadjcYV5ApCu
O41zSkOQoH3vWHidreePwn6sooUigjGP5zPi/8YiL9GqYWP1bJXDaxAG16LtUVVZsZrjR2UDiARr
YnOMLVpMJUzU8TzPwy2hEXCznRgS6/0sDGrIZxiMfbL2/omPpaO9J0mgD8qaly8R+T3U1Xi4KWV5
9lCk2tgCXtAmFYugkgOZTj7LpMFSDvl+XLywUrQkYk3mdWKhumcSsRHIp4krHXESTl2qscE05pf6
wBv0UKbcuzDn0+erOvqlenbs4hIuZA5XoAEuKiE6Eipa9lwrUAG3nMMfeasC/3ZO0lwN42Xmj/hg
xgZnvCpTAg9V7bYjr71C2pC/YNNkE+wCyUHDX9V5vzEmKUOpM4NmuaIb5ZdWtwJnrJIGLRAd24aB
bBOaHAplkmXtfcKrt6TwEu/iQRo8G/t5vWQJJ3TKk53J9yooiiJEnvQrUTF+y56dxjVp/DE4meAI
oXIfAjw66t6+nwyd7kdO6eZuQrhrvaqzoVGdJR4EiQoaBQel/pVNCT9WC1zg9urBmpnJGXT1kbyH
4n/fptN/zlgSN9FIVQYFZoh5cn7Yi/smwryf9RnRrWafadx8K+19L+qT9gRA7aNnYirgznN6PNZ1
DtRkPv0IzCcs7b7zZUtsK6I/F8PuZlKsRwfOshc7KaLeA3D+eXw5XAjg/fyOX4S3sS5W1Zy4ML0h
s2Jtw1/HTyZ0CylEKhNc+FHfhynhpun9FcgEDDzrUbavpLyHotdwL2+U7dJGUQXuwomQMdjkH97n
5EUY3CzDaODoPLsWXU3ELyBlPgavpJxwyRgu0sSiIK3TT2v8uC7JGxh1BSPFJsKf4nweesxTkagF
0H876F6IpjWlxZT2nGq4reTD+uKfTJ76ldcRgxAZ20ymgwUIq4v+cT7kpCqZbK720JmE4F7X4/YT
q4eEGa+1NiKSOxFtZrKnYane/P4Hpi1HdLBvMM14Sxm3SlyBCbadcSfWEJirnQbnxLovL0rW+/yv
HhCDC7+p2G4S4DBGMXglZ8LG9ya01XmlvInWenTrLbGKS9lBGy3+oi+VYJdD26YQd9Ff9TGWla2Z
8zAUL5IxpB0DeBIvhwQXKF+3lTCvJIQrvl4FXCi4yZI7zCL7DBobl6g1UGorRPrOyKC94jM1DjeA
3wgu5KhA5RIQMv66Fn9XRYIo9DXNdS2Le19SwItiQHj5zuPyt9EBJk5TET3g/raxUr6DFs/Bqabs
1MTjIMtnB6I1qjxmCvGtKCAlJBfdiJbrHsWZ18cpL2ZduYDugLqU7MIYvyykexSIbWDQWddSeMch
eLW+Q/UEdCgYEco59msNLEHOGRUhXbbdScSFsjpcT58oUTI7fIBxrxaIffk4SC2VXJuu6icd92m1
4/79ihYG4lG9psoJUKIglqdkyX28q9lL6G4AJzWhEw61TNxcSCxPAb2gc9ntmCScMfNcKSU8Lj9A
dM1+YEMNK7VJPHd6xSgoODtDsebXSWUI3bf+/vud9++jPVVl+0odthfOGd6IGAMheuTNg9F+ox6R
vrL5y2Cg/PhiNtLKz5Lhqucl4uIcJg6MhL6FPpY+eDRo9+CnDE9S0hlXvkzhR/S+FpjYQxtIST2x
3ci5l8EMuJuqNl6WGO3ICRGtWIo02LVD6v63J8j02DZrAHmGKKzT9TQZD+sdNxUs4/cyTEQW2w0O
C0sEfCEsh/3A3Q8jlJAkWjQ6KpjMWQkp0cUemznJbNqMrAsTGHyDxLsTM70pwNDuIvtOJjfQWzdW
jSP8XTgiQSM3l94Kho9G69K3tUmGUKygUJkEMZMeBAE9oX1FjuLjzV7ac24lN2hlrGR5BH8Iv2vN
sPmLd12oLx69yXAi8CGtIM/R1O9Cx6oh1vhgR7tv41xBSlwmvk77PEXH8N6MrPZe5PY86yJ05A2i
K7kIdRnaw6ly+j1LWMKnR9gYcwD1lHqHg4s0gSArJ4lyI6JCoqLK8QXR1bUqhvhZXNJTFW/1NSE/
Hww91mesfKHWdGIEOXh9MmlW+R9Nk3Xjax2JtSThREsLwZxoSdQrzj1uAmJGsh9Rrb5z7MsM0i3y
YIdwYnONw/1UF91mZ8mVgMlFZV/jHy9La3IuwfM1MpkQIFQH5WYnQDtRUJ/JjFIoOtM0vTizS3rq
KQDwlAMfIv1H2CTiOU18B3bwuMyidqqFnKDe87Qz2vXGxfBq6w/57WVW+YQ7jFYQ7wKsWnL+MsEx
MihOA+x74Bw1OeQ1OZ8NTkDlAXuVDCo04i8W4N0wEBFunwwHAJLFb6kSapHNohsi04rgzZLBTDMM
YIXrj24pUPVR0lJvaQ/WhdsjQFIZT8hSF+q7nGVy8KvTUhX7qQ+uo+GZDQxDhNupwMvJOzT3M8c1
5eOkshgqamVOZ4/ZzXqe3ZTZRxx51MONjvv8wnZN3xlRAryDHPPymlDxErrDXOGmZau+Chjw+d5Q
XhoCsXnK9J4fSUXGuOuJSEh2/N/yaWHATt7D0h+KHAnkIhYi+hOhT4mmrJ/D+Y2yO8nV1gHUAaE0
Xw54SAjJrwhIYORKhL7JeotYOCRTxWLhx1WP03gNFTyGJnDnFjIs0YzwAi+/LvPSNXPsecrDX5NS
oXl1qyFnmInu1TUPVznMamulySiDUPoj2IriMIlmKKOwqYzZG7GWm6QeZKt+90ISJp7r9xSwJbCd
+WIPdJcjlSAnx2KHrwRBBZm6PAv7O+MB8UIx7LXZq3OM69Uvwe6FUtlSYXTzfTEg6ucI189gE58K
TnUT1CWzVvFYZAW7uxeefMbnhFqvJNZSIfzoM/VVYbRAMcY26InkJ7s1yj1JWCGX1LOW5LcnCk1o
gMUrOk63gU77GXGAZqQKoxUJ7VhbgBEGTcgsAvuU0Yu8Srk/dwLIas+cJTkBi947JeiMWsJQv0eH
kAS42egDevTJXtNA6zoU0QgLTQyvb5uZ1A61Evtdmy+nwNH4IcfLpEw5cac/EXbgCCtXKxHoF5vi
SLj818hLOuBnRE18JDOKpjPRoYBxVpO/1mT13dy82YPS9shBIstlWBGUWFiwJ9bFjewDznMc83iS
gVMwQnrUYB+GeLMpeKMwdDe5sU9LBCsjKU23JQeGXPbZ6F2+cBNfYzLe+JfiMh5BzSpUZf5jYFQa
rJCM0TeuRPaFmDNcrAo5bIqeQ4T+2qUuR5p3+tgho7K5OFEVrQwzrurH7vhhwE0NvhnWj++iWp1J
QgaHRJX9BdYwwmo2ILHiNyjBNYC0jsCF2TuZS/oeY6xMVI7QI70pREbrlNh1DRF9Co/ltcfF4SXB
IH4n0ADFT1bQBHr3zWUmD8MY64bjfQ9D7zKq38RIeTBnuNGzYe0Bf1DAvV5CADO7kZTCp4B0ck+h
KgB0YWZMk2nwMy6uOocBJkq6w1chBtrGP9d/kiC+e2RWHlKbcwEADBFRFn3ekZ8eBuPvMpA74eF+
RQskRhzZqx0cz6iyq48UffkaSJbcb60rCYKi1taTSFCe6/iQYCypEAM5wV9nXA5AufF49edn6H4g
9V5+Hu4Ndcka2ToZWoahE6SjQujUX/w2DG+sPGtXIwkZfGxWr+91z+ooZETxWlY4MfzctyXov5ma
s1yoMhfhPaeIp6hWPrJWQCyABZqXlrufflQBKifU0Gj8lWqInis9cu1LkHcZ2VVNILVA8PbmBy3R
6gXoowft8RLBMWRxHxbYAL4EkXmrjlxcEvAsCpNBNVRcPMvpFatg6NgL0WG+9jgWZbmlRkBwM8I6
aGQMLjCldDqhB+zy0RzXIGCLy2enktNnMdBrUnlI5MaHTNtGAhehUdGsj2cNkMO9et5uuQKqr0nG
hV9H+WKK9awwDMZdIlm9/a4qYqVmSacWNUkaMGMqRHobG3Sc0ArgbKq9bZLCFsRUGysbsXb9x3IV
RK+31mMRxaOgdMtScV+EvH9WQQ+pSfWoh8raDMW3sFONKN3PpQG0PMdyhrEH/EYJhzco0tf6gdLF
KpeuNXqrc/JfucnsBceNkTUgPE69N5WUc/NDmYlRSaylFgf08+qLB8A00l+b4vvVoS37GQvsXwIO
X5GolFvaViQVF6IJV5lsQIQce9q3mieC9qm3Lb0DMSafAt/js5GR568tliaomu936yaDteRG2ZYv
PZSqKcdD1L93VO2fLFu/VeRPmQc8/9Qq+4yoamORXIXXFy7Shm14PFhQ/xcyhpk1WFsTTxXrkxvj
z+8vDy6vv060BO9SeACXpqX1nRnkwUGLfNqRvmjsAdMJqwOCT77mwpqUVQIaWRnwaJDKv0+eMTw8
G9V38Thuxj1u8SV+BXwD5IA+qGV/d0VlGpauLd9ZafXWal0Od6NuvY+I3GsAawZu+Rctg1bRKKPD
es99qNhVHvTXXcay5bI4fwDZRa1Z5xAf/8j2HmCAZcTs/ajcUsV+lR+Qa2nzT63Nvb7JP6dWi4ek
Or0zYU2ztUa1EUqtwNM9RI/vy619LGX6dHLPcvJo+kGYbIqf7IoPDNrjNE7fFqFQI1lv/spcPL6G
MEbTxTEvrMJM4/IhMSIsyl+pWSL4aB+VqdV0tYrkywjNeBlMMu7Nun9qKWy/ampl0szaTwie+/Ak
uPXVM5onATP91v+o6oGCH8fFcTKqGeWCEfRmgIsbCPkvI3HTTZHQ/3G2vYzXSAsS1Q52Ff0w9D4G
855PhrFxEATKeZAvYPNLbnHdvURDFZDZW0sazq1MCmILQlrkh4Sx7cGnf6KGhRGBLUgtRigkV8L4
G9gSfrLGOObh80PNw5G73PwHqFhn7hAhpWpUgSlewHvdak8acpegndkHoG2O2wGifSZbH7ZrwM/0
fNYM75kzHR6AG04MQ129ibCFFmUBteFP/gzLlWDtm8gWFMGYQguCcF/ufzng3Sm6w7jRBEGKUTD8
qgQaihq7XvL3yhzVdjGjjwO/FBnfV5FjZh7pEFZ+DJhztPaAJELu/xBME65d0WTz2SAKgVIfnwik
u83tFC4/hRQnZYaK4VvL5FpSuHmfmA3tXJS0ZB9/2z9gVtWn+EOiOOG9fQIOpn9spMqEBREB/JXg
mHhJLESG5bmd1h6rbX7SDALs6XPvOQH3vb2+E0tn6KUAbYiPS25pKfNRnsoQqp0SczyiI+8q+Yjk
JW6qO0t6QwmJ0KN/65cJG3GUeSHA9muu+XsLxZOywHeiiFfbOxe5ON5fkvXzkkXunthhQeH4HRyZ
j29kbAMaX2XiXj4nQ8dH0S+YWmt1iXR9Ek0s1UnAS5Fi01EgU5/oTLFNynSLvd68JhVK1YQWYwJM
ISvnzOf1AHTILEvwJmIJmMcoBzYgURgiP4zYZdIisDPpYLIIRGdsT+8bN2imBQVhn4Mdc9WWrfY/
h576knBef8U2TvTXFZhJKcsQIEsZ5LzgUDrTouq404ooTUsx6MQkIXq6UF7ZHsUznpAUb67JFxuu
5ka1aU+y7aRRqHeWX7Vgp9pXisSXd/L76ZP+NSSI4O88m4MXsYeHs1Qpj3CgL4bAhXr2tPAYJNNd
PxJjw6xuRo0bOmRgdmIFBWwhjZkrj7GAkONdC9NuzwBsVB/8YeIZ9bA+QSyvAxKDt+0BPCkf2euC
/4iCyiUvugD8nCp3r4OdyjvYphw/yH6dgRjeh9CXppC4UPBTHr19lJ/yhdCJ1CqJlLGjp2Mu5RZo
f9lJPbr2s85lfSLP2GDK6G3d0cThos6nHX1QnM5jq7+Pf/F2Px59KG/GtuLFJerjoG5+MouLiNwj
9z39IyeT+SuEyHA/Zwo81yX3hPgzYdaTpTvNgpUDv6HLY/T+S4g6xAsaAicLz1+iuG6nWt1rbRgg
Y41uOpsD/S52GbZa27uLjFzrSLGaKusWYdrBxtrQ+60POQyIHq8lXTO2N/TTF9ss0a20HCf7eEGl
vcV27yVN9tG2Gk+YoOULYeCN8xcUXKWmnDtKQwCrDHF+SmkJ2LbeayMWXE/oNCPDVX+DbtnAwTs5
DoJo4W++7kJOldV+aogKGEOHBUCg4jYBdMDjOW17kQnlG+vegaBqvJ/yZBzUyGdVgMYHBDbPnJWp
6uHeFvl0BRr19crx5WI3UVGmbIcwM5BmU+W9+l4aRxI4w3Cpzn9qe1EPRA24AEfhjnpI2A+hQskb
o80bFkwSZidSwmodmq+BE997LrxEPZ+5hHP6XAZ7oVGha3S3AFE0a9/NDG9NQKWNyHEwtxxRXXme
+t53bIUAzkzoYOF9vna/x6eMAfWndJzhsCg+G2Ke9S68QfGkwzgbVkAhmBkeU3xykM1jutwC5+lC
UzH21mlBKT4Pg2B0W3jSRklm0XY1fM/x1PW0CrsJb8yLSMrVq9KT2Xuk0NyyfzupiwEKCDZipdPE
2mH9+w9XPuv/de4u2WcuMzo/zlLQFTPf9SyrrkH5+f/2pvGlGDY77BszNu/P3iEFZzpLd2IXj10v
ZnHCZF8U+GirtwPzR4fxUBmEwQiwHJN6cQBpxUsW1D93Xg+CdhuYWm/bgZx/zKCcNN9ROYN8DqwG
nePjLhIcATJl9QTRK6krO21QKZRSZ14DDTfTQV9/XqaywrG62ZuY5wDzWsywH3ERSAgkvJ/ttOAk
1L1SyGLf47J8pklyHNgz0I+R06L/O29jU7SYxRzUtIdwYHaxA/e/DCHK4XCzypnJUMD53XbYwiGi
6osnzhF9thd3UJGn+srbRRqcXaeaVAbTNulblSjeR5QbuhSTinXKuxRbnexYAVMR4x/pJk55KCwM
dEg7vW0/zbE8DR9l6KF+7kZZn67PmUsZr6ds/fVz5osD2+YLQ0B0XP8n3l4ZtuCVf/QK0guSmAro
Gl4ExqdoGupWg7gCB6NlDIkVw2zpdFPk/t1pmi0NAtDzr7JHGy/CCco0nKbmRQ0uXBBd/UoGw7ok
W3FfriOyRwqZZvyOkEQvSOaNMenJ7BQ65QO3x6zeGOGlMrdnOA7qTJsfaafGvrlo5gxyxHnS/2go
ap5teu3uVi+qOVOVSzW1GO27o/W8+awAy+pbjeDXeRGSyMAhwXl7qPULmj7mXmMerhadqNBc+Esc
tKdo/lr6v/gPo5dOoKiMi4qFVqAaTkVr9VnAULpvvVNVrdhpTxHDi86Wkv061VMIwOviWAjHw0nA
7ONiUkyyFUdeJrkAOF/vnU/bU8wo45DmkV6rEYxLmrWr6srjUU6cZSW2XqsQLuB5/5VtkHNIjhTL
lnHyU6MZ/H7blLr8oIc8/J/R5QAOgVUat2fdiMz6IQggaE5gsSfSJaExJgFtC7L/Dj//NodtJyz0
yvhSHmGCnkoa8yzZuGe8kmNeLjTvEfSSSGNz1TOLjhv/f7dt/3j/NVbGkA+j5Y6BE2HKQd4+SyKu
HSx1BF5xSPnQSAgzRS1aRKvN8PA1pHXyx698b1e6whiklcoqPq78CoAbsmEvRG4ZOCOnnRtFpHhn
AgWcalVGklKrMUtUwz/Oe6ZK5uSFVbQDGPvNu7laEbxCFB/zFF3bw6Sgln2anFmfILLrB20pujfe
WK+DufpdrabJ5xpnuylhOCVWitxKbKIJH0AS69g+UKb6yFUfGp9vvVA+GcYIfcjqWJOdSDz5D9mT
c/SJjq6RWYAn59FdQI0cTBXR0ovggPHpG0UqrLxBx1X2xY6SL8FLDTFL/Fqh7puCKEBHwrgzUT8t
HPv6Ox2M6OU3iBGua2l2klgsTvRHMDUF9tm5ngRvgj3AlmsJ+ekXexDzGKSEbCjDA+8ayhqtCiR4
eIew3JxZ8QTOK+EtUONfRkkYNTfvCQjLJyTfOzLK5zM3YV0qrPozBVFKSMNR4iez4hN7NtHsDrmz
1MUqXIDLglSFegpAt4vmfVagCfDeRUloQwlhS0d4Z0PzAq5K+FlTCYqEQ8JSo5YBN+VzvW/aQjji
FA5Wk3yp9QLB3UzhuByKtI+vQtQgW8ExlC7NbT3q6hiDF6cIcnkC5fuZFWT5C53WilNjTnklCKAT
RVZhXvxEvue5uB3MmseVnjfGDx9hxnJ8TdMKeEDJR7rJ0+M/Ueio0QTCVKF2fHQcUYMUX7tTa0Pq
+hNmstV5nzdaXx00GdUdmJsv34ouPQhpZVfCHKPkeODkkemPVi2p6zHYWPLp2n+STceIhsQSrS22
GJHMzusLnT6Ih/1lqSa6lPFIbxeNOeRLnN0scchwSfuHGaJfM5SZF/mmCHggTf+BeWZ+xNnj2uCo
aKNNOK4ARvxCan9jsktpbNHzPj3B+j9856bLTmVpH9f+xXS2Z76aRe+OnX/il5YppxtGLQgsQ58r
+C4BayCDJdue3L/o3u9YW+a5r0UaFgixpmxNvga5pQ2Uqkn4uG/y0DWQlSFsEXcM1YPEaSx7jegK
0sEzInJr6WBbgX659+BjkWOx1+IaQRxT31nPpEKuq9YyW9NpRPvK+KiHmRYPMmuPltmz3wdjH08I
leppYMq2/DtvF0w8k0vQQGn90LAma9B6tO9wooOucoEs0qvIZoi0YhC/J5c4mVklM2B2tAXfVW9R
pREzSWVaaFTLBj0x1uRlNEOmZetwBVmJV77SfW4TtEF3C6QsdthWqhti1pVamzugsJvs7YJygJSd
49XYfh1MGKZWo595M+/YZmbnu2/S8hFjiWvoDWNWSk0bS5ntn71jb2YroaPrE/f4ETMfBwtUvvW1
bm3V6ZIPVs1UxcdWn+Ca0NdCChQ8gSZD54Gxz7bYC7hK9kf0t2JFRUOo6uCqfnu7etVYEWz7W1bo
vSOjoHv4XBvyReXfrxI2b5QLa4H93f6vQ6oRjofJG1bM3CJ58xIo5p0AOJDc6+Fnk3ISuMmDJSaE
guC98iSFfdJvdoShZ7nd5Z2OAWm17drcfW9haZE3izBZ7p/PtJk8CdhhazCviXHVH/oHAlkW8pOX
TwDt8537eecEEHbrJAa1LJzMfpaKqrMoeBNrcnLOQ8cBqkb+xxhPThuj5ftVyEZK0iJ4juqmPEuA
CBDq/4aOc6QGHS/EbKHSFKep/m25lrVSV2uk2TcYwDNWS92riHoaokn+HnYPgnIzkadM/DS9tiJG
3YfZ8lam33kEBy8+jVfIN6+p4X2OA9CGQ7vYMLcEHYXEcwwdl03lKw8wk/eSllbDwjxWtRLp1qi4
VqA2zAR890X1B42njdBw0KRmf5g41f4zOVtOoMWSHO4UAbnIgs2cyaGAqgH8lVsGclEQPvoykVjW
Bq+mNKrnWF539LHSUimJuOjDXockV4o1FfVqYJWjeYOui2yK6J+tskLklZkFebJfEVvmhim72vNP
CiG0aFD3uciVI0EmUBbUld1jZbXwRkQ84jsO0p9IKDBKf5zDybz1vDNsPfWxO/UrXUAnRvSYHb6I
bhTUlh2cPB6wkPukSemHNg9RUfygxDSJ24/29MHoK0h4WOGGZZ8oYP1bRus+yiUNP1XOpC1O7zpZ
nSCTYxGYkwlyL9AsfkVCerdqQsRM70u5+0a4YSI0Xm1LnS+IweLRDx5jSNOntZjZsfxH6Ps33TEr
Xsyx3QRn4ODak/tYNjEx74KZubgIqR9xEXI1m0Z9FoVIkkZ0h+y95ZP2igTPO58e4Da2rTIfWHYO
NkA325LjBlvJWj/14mLT5DcDKQQcph50R16NnVFQGLANhos4IaovTbCOAOhfkv/0Xf/OWdh7t81t
bK51und3QJf+9braHmw5jTTGIM7YFO3OPpZzguTEOLzfA9eVBK7jeYUbYmLoyKi6C442/wYZUkF7
DBM+BAfvReHUYXarFZD+O4b+yAuGPeEBYq7Aa0v4q/4nlq/yClN3MnqlTRgPGT79thZSyPwwYZ24
BHZVifXrahtKPqT8hN2uOIv7+lpljd9KBn/GWs+oSkt759lkcG5+3Ts6ETrbi9GUM7KUxmUOKvN4
yys41DPFOhGDQvolFI3P42/yowr/07vebD0qM3Rbm2kgZoLF3qkjO/Tf6kfiwGOxTwllbmG+7ARv
OtSO7QpP6xs0eL9rHUrPizdjq7r4Lf8YB82h2N5j9hwVXrtv81wG0WQrGGyJtkeQiQnti3fJliYG
UHZG5Q1fOrCJwXvB5ysDpv5KzvOQ5ogv38hgcvDcH/6XXbiRqoeUzFmq55eBG76Y2ydZCYEGMNTw
msLximxlbwaQ+cPcLjGevYwBJoaeO71CQLLVUz0Hz2Wsgsn8tRIlAhAcA9Eq64m8EFN4xQKIdtrk
0kGI1L7ThUY5CgrAh1mN3WjM0hD2ijh/q2Fb9u+8FTHaeyvzD/fjTr3l93TQOD3/8eS/OngtiUp6
RCEbzyEbgLn1rkW815dRL2YnpXgT9wQT1IAq4ZWXQYog5caUL4mIeXJhB10AULmp0mI8vMWoVBxe
LZ/0j33UrrhG5g+d+W13oCAIveTvl89tM8zAo+Yf/XgfCoXWZNe1TLqKg2wCuTReF6pSuDRC7hYz
Lz3Zo1qnBPkyE4s0LpbzciWttXBjqdwplZR4gIrm9m9kt2A69fEMUciVhv2UWHMHeZi+p0lwo+bQ
S9aGss/rbNypLpKQBWoKUJg2oO9phHv9TswkSeSM8jN56wTxz2xBP1q14Y3N+iVmtgCrTtc4v0jU
bqwCYHiRjlpdHbHM9P9jJYKG4Y8QNKfAqSLmzWSEAu3ii4cANV02M+mVDDbWh9VV2aSu+9phW7O+
c8oA9tEd4aIgXp93i++XZxySuCJerr/aAKGTPw8djnns8kO7y7RggokxygMUV6XuKXDDqWgX6MoA
C5ejho1t7SXc3kbhKsOKHh/I8/hxgepXG0jEv4/ACuuZxHPvCxV6mm2VjcfI0HAQZOzMNHfNFkH0
NiDQERYZygp8oP6WAgiWQdYw/hYuXp7TLl+jkAYXyQC4c9A2UPwKnjP5IzUYoPOKDTf+vdNHj20z
/mOAtETCVVs2Ntbo2rny14xZW1tEVuZOK1xowfxjgYS7cjoaUOMjSWc79xwwLhKJ1vmuBceW8CqJ
IcDto2xpMfJ5wpteExU9qx4UDJOJRDzWBG6+JS70PHE16bicpmvtMFWy8Ug5GR1YfxJnhszlV3Is
gWdaYgyr79JPi6KIO8Kdrdoo+Jxz6F4ZFBsz6LpWGOSoel3ozsySvlceNL/rbM+Xq+6tQ+asSE33
z4EIdVFuIDzzwJd7bZTeSDs/rLPXd2hrU2a3DkgtqkIq73fbL+by9QPNyKkBive2QkRyC2HrAiBN
tW9r/59uztAlCbeY16B7tApYGcc+lol0PW62LIus1seyH0xtanunvF1lQrqqGlXAC6uqNE+8KOIm
nMxTGKrSYMMv9NBrZ5L4143MdXqJSYqx2qSp7zgQijr4mhzWI9dPM4PfPhSSYrDnQi7E3S9AzAD8
cy4zfmvYNKq8QCuuA4VR7GLEaMymr82SuI1xWYFDLciyYedDcYQmR8baXbLCTylg+qwG+2I3dzif
MOeROV4KdXBsFIR+wQCgMEiI69fKibDBeSVlzakGJCdR2HTWM5VNrUEFXx6yOFu5KJUNFLoVIZyY
snaPKST11W55BP1Jo8ig4wXxR81V7kL/QXoTcXWeu129zd15B1u27wWmMmcIxuGQhlQ0gKTGy5B6
JCqyuf2DK0ORMaI078p5VzVmK3WVZiVbZI4STBltrNTRXTDHjeMUkw6PwGE7CKWDOEn3wyy91QLS
KSgR1D/KxTfgMNBHwu9dF0hOUKjfSpnNiWpZKE8Cui3A3lyGP9yUZ2g2ORKCZFzFaQTWLCXJmge0
RSDNIKNvPfcgm1Llm6bSpatx7foxZ9jckdDBJACuN9w+iPrYs/ABsp1wzeJU49n6qAuP2gKtRXLg
6l23acv581MQyqg2Nezv62Xqt+r/87EssN4BqS3pXHnCmaeIoSKTcfHXi9mx8RKaisb7uZ/bbxIS
XxVS9VQoH5tP81MdXXwOtvhdrrmxAxn0sBQJPphDRqGnrMwTKAomqi1NTNHOHINl5H/j/AoMsSKu
o+vdNUuVN6RozJp+59F9tvqbGhC7bZ3zvS4nziSAPgUF5Rui2hYGmdjZtE1dj6fx/mcO+g5ybjX5
yOvMEEQSYm3uHwAklN8TjAtmr8gKRcujwMnaLd9EMPCafVLA8E6JIb6G05pwZx8o+7WHokL3xvQb
64mHzhndZzzWl+noiZKLdmtfPbH34oNpdQ4Zwc8ZFLRvSzP2aSarjiT8I2/zHolDPMIzO0GBjW9S
z2cQHKa4kGoArFBy932SlThGCGpSWArvgfSS2XsZesfMje3/58wFoGB0PsjjF7jaeA7jPeplgntX
9u6ew76ZOKP8M3iPWbmemtOmMnEcmEYsvKo1FwoHO8Vd8mey7lKguyqJaDM7SbtJVkxHpAHj1gLa
TvJtIwQkbOSOyMRZTnl8LgRVmHstzxpcOkOaO8/ukubeLLvHUhCvXN/Vp6Df6HUwQXEbTSiYeGA1
oOQ6MASFmexGnuWJ5g8wjrmWqyucsE+OGupKJhdUPPUeYjTDwl+jB7j2TFsc13Z9z19aB8u/s2+R
0TAV+kWM1XvpK8I/ACudQ4w0hXXDcI8Um8Qfn/wA+Rs6drF6HZTbEwHurEv+anJ/VzqUcth0+nwZ
S13yIup28iIcqM8sB9NZTINzmyc0lxF6fi5qqbUW8sOT3KEZAd7+yQtCAue4y2SDdNgd+n++6jS5
/mRzYv4kvKQjHOLbsHuQK9ogRwjuH6DWWjZJpYpQ0ndPj7J0GhhE5s46qmgdRsDAoTYfP4Sibxyt
HarhAGLjySAlcs6QENqyx0/FpQATKXBwttZiYU3gTAZ/6uBl//XRLjqeBm/VviD5TEUi7Q+QXG/1
kbyA9Bgh/V1WYUyga2JaLKM12TXxZszERb0on6VcNhM7I+6pLe88/Pg2Io/HetMrorJa5Lu3L4/S
H+3yt4P2QACUvZGqcGT+K8AnYqh8UbBC4KgyN1FnuzcfamTgShala6v4FLSILqWfOcKmewazKUBf
tYXyF9cKoIjo16jAu7ilW9izmLVO2L5XaRYi9X2oNp4B9R1Nv1q8m860s0Cm8gGOagUDfSAQrcts
fSF058Ru/N4DvRsTuv2eGim2Cehc3dmieRbSV1YpDHb6aV8AcJpQ2o5QvAUdkVnnKiaSFPlBmGU2
ex046G8X/Zv3daaz8fhhsUkSNtRMJGQmsV1A7UjWYZqK3vKKRVKRvqFOCWcMJhu3C5fI3KFjZEhi
yqelyEdsdGUq6xMRXkLCYEVExjh36OMVCFONXyWSgMT5sCkGxO7mfnuVaJhSa14WA3pTKtFvh+0a
D2X20VwOSJ8BllDsfjEGJIJADvNObYzhwQ5KLH0NLku6PmguLwpLdIk8dUeNPI57J1u7uzBXsK53
4pzrYNYByTjrHz3oybwJAg9OeJJvVsG8zWEJaO+6vZCguG5Jw4fgPsU9Mm/bEIUAQ+2q+y2KLPqk
WUq5qBs+sz0T2yBSIggYIra16oYIktIMK0ZlOuQkaNdHul4ZurPQCS5GfiQyWpxuvqlTyXEj86ao
vHUvw+dwo+UaW89ksNEI1e12LlSXfAEKkIrkS2zEGysQaTMQhtGlip4mYdVAIgp05+GpwqUHPpqq
TnWwsdm5S4hryaZM4Ec2gyLEZodMRxnEaQ/oeWIwUVhT5PWTdXGjGBbmfFGPlN73dMdFSiBxxfRq
JVQ+GHzkiHil1d4b5S7RMRzkNf5QpjWYOOCAJAWWuirSK8WIh+TSVpWaDGVgF0C40/pconWiCros
zyZ3eP36EA8agpQhLAehIDGx4m3Nv7M1HD+6KWuRf+SjaBJ1za//gEe2Ji863EFdiWJPH6lEK2dk
8NROqA2G6jnhwg21eUlLlh34GHKCVrQoGH/VwbayYJFeReoE2Gq4QbxmsNOuuGQ2BNi/PY7rCwmk
RdNQRG72f5fPF2CzsmAXboWp/mRvo6J0Xpm7NnoBw1VhPmdkeu1IZsrqkpWBGRXU9NwmL3tfZEXL
2JjbQ8Joc/M6iymbui999sq8OztK7U9ILQ5dgIrkKVGa6R+KPJaiRtgGPDN/6/rJltuUDC3qycQs
g3Q926OKQdyZYKRThOMJbXfOY5dKy9La9q5Fx7xnl8pcPml6qMmmsfbB6m3eQvDXf8DnXruWcYeR
QPBApoZw0+XpLCST+SrBrmkpPO1MvveciZVNk+cRRHvXQjCm1Oht1GecICRy36PyFetSAmN9+ywn
s2EzSWDXhztlIRU6ol57XqZe2VQbLpmLQQfHZsWTzPik8QUp/B6DhFBTJi13qZZlyt+34BkNMiQ3
sO3bHHLXMGM+X5faUQ4lYr9VocCNhyp5PAsjjs2rxmVeh73ozfKubaW/zNd2TYL2tDyXpLJikdqI
h/u6brcEWfYC0Xgd73YL3gCXuBdBoPc6zGnD/9MKh3fy/gfX1FUN5svn+dgpqPQs0wbHOZc9XvqU
DdNhxNuT1gwptuOUJud90nlZZw4XWZw6jjgbwGIXe9klY7h9lqJyh8tyrDrjcviBj8VRu9vl7mUY
PsVgANrcqbokBx3N4iyecZsCMURTl+Q0i6DMXgIQzHSVA0VQXTHCAIKeaf/RzkzYBrK8RYyq9P0t
G6dao9q88WImQ5zWdG1coCsjs623R697UwEerhEmTq1dnLA601uXiGs7YWHc7rXRLwD6znrAzeKS
/C+DM6AjPl5znYNiIDfAjNj4AmBnleKJI4padE8CVrCc0LBMXzTOdo/iXVuMtHptTkHCPnpTUyJs
fIJoQZsEuXIAtsCOmtbHVSOLN6ozpz3ad4WY+ND+rYDK/gn0vgKNnQlNwM/RNqCc7S9sgd/U/nsz
xsd0W/nMR/WvYgrG8iqQLtdCXBBFaEf1NeX8nusjoWtltftsxRoOymLYcEzcd7NXDjrfOkxePHKU
SsqR7mpW1CZBnGw+V08ZkmQkGH/XcW5spXj9Tog+4QnpkJc/oKtOEJ9ePsR68DSDo3GpaiAOg9r2
0gxJ80N7OmMvDNHQonmDVllBqg1cRItCUwd3jYwf+s1TKnCC4tzFn40GJneQ3Jzgq1O6WIPn5KQ/
b6B06W6KzFvSw9szVmi/ZpXg6XXTaggH1cVBK9G5DHqfUWKLyD1ScoTBtXYhDhvjW1YdZeHV91R8
I6nWWHM4G5crD07ccyeu0YjwluEDOrGAU05XuFCnrwFqitLVJElYsuWwUIUpDG+5gDvjOyw79yCy
ugEHqXe3Wc34R2xAqjnT0NGSA3Gmp2CkLFgzFLYaKj6jPJEkOI8QJ6v6yDs9+0y2hnYqYNQfA9iy
+6rvJYPN6G2EYbdcLO+3gFDDqmD9nybPBseylPR6qRCqbfYCg7Lo8pEaf045nPsnmQzmOeQfaDQ+
u8Vourufffnl3AskMH0+aEKn7jaRsIA7v44rhtxdmZrwGrm7Wu5v3VaQNAJXM1XZFdVX/fvS95Fx
i23H1BZlLy50kIyR/BWYRPfxHPJ6+ZcLut2hvZTV0XtNH/SMhn1L2qBnxQhl6YaMzI39pTUBeFXg
5c4vA8E71vDgg8LmVSnROiMeybXO9gd+PxoLEZy4MBCeaaQhRtt2D81ckVuV3mj/rMPJCpdzKg1I
ztKCdu7solUPu1e7MjLh48DW6HXvix+FEj7pwCTFFutyZCi7FwiePld7gTdP7VXGjr4AuT1zOnKw
5SsZQsmeQXBue9lOT+PHHivDdSYyrAyyvwwN1w7JlswBbmrS6R3/Oqm38Q3GWC8A90th6NZwfgNt
Z3w8WzMhZxoYmGNzrSSMiwtbBkNgpkY+phpO1Sd6fBNrfGNhrruzYCCfRCWGQHeicCgUWV/rMKMH
vRZRdalYTRfVzo3nChFFMO4zaTeZ4SgCCHlBdGD4vfY6e7agf9Wmo8Ex2QhMBIAz0weeL36MyP0b
suQ+JGALsi9HdrG0GNTWBUNsAkrOLdJ0fsncQKdSgT8AqpAq7ysDababVWwBNe65Oq6B6SzQzvjA
vNl7aBIboa6i8VjLp0hZrd5y+1bEOgeYA4iGYWQVDqwM8H1zcgsTJ3w2GnvinRwd2VPF3/xIztE2
1p+78aNjnh6YeYTtjzVw+OdT/wbhSX4MqhiK0aWYI9ir7wyBWHE8uwepvWxwywNaTiEW8eDa/WA3
qINDoL4W3XjMdytWeoztiHua++mgzjnA9lKuugW/9SEefH4708BHVnSF34MasWm/Q3YfMEIGycuZ
IZaeBRhUbEVm8zATks5DTcXfkXZpsKeGF5yyTgpWbfvBVen26QPdevLrSH6kOj0o/d6LFIUn/vlM
hHw8zOHtKbvFUyrN9L20m9wKJAFHLIyjOOph/69DBTbycbjcJdWxLlThMicGA8jTd0Ym5pe1Ak7t
xxDHvzpfot+/x7AROI9FCucDvWvvVOUkUzV78OSIRX/jVm4fNMbkai97bY7GERfnTgD1Aw5w7NEL
io1XE5neDpIBYyOkhxhb84uZgSnrtEiMnoxYKEjPGPPFXiKbmww+ImeJNdNl8dU5E6+DpCV1Gy+U
dhSErglNJzpkbZ+Y+VYeagG3zFnBSEKgiOC6nxsMcuufbMvJKOxzUlSa6zMCr6vyFyYt/QJ/Q7R4
bQ/bWjx3pW+n0CC+xVlbcXAEaQlOfQQ3BznQOIctzVPgH0JELn+Q6Uy9e0lbo+2G4SjDPj39TYCv
BFaWSrUT7en/VPCDdp04fW+uSnTuLhXBMOxvNV6wecDAyI1C/c4EbFrbI76Q5nWwGj2xC4I0wi4M
jptwxYxmFtVZ1rqR59qnQwPaV/lgyzb4ELdD7gFhUAGNVJpnGMTFix3C/YzlofLvLAB6DjpmSTEB
o74uRNux/o2a+eFIu/wqLIEhOZSGh4bcU4ZY1REVnUv4AJhXQpHHLpC3MTrqjo7gKwPLUFntbCPp
ZEL7h7uWvbjzQ6NaOeqvj9FztoOVzJU82YW/oHNnITCT9cVEkXtrkjJreUYoBQiQYHGuSbxpaoWL
QSn7Hh1P7YqDAmev5LrHe6hZTULZuVHeK/N5+W8xp2nfHrYJtvi7FUnhNeI5CXimdt33YScD7V5o
Mnhh7sE3SwF22I40XNBSPx7PCiljnWuSzYExHTf6V/dGs5x6dPhkph3+Q8MFSy0Gc98CYq8v3LDS
+I+mOeAmNVo2rCaS0crEYjp2shg3mK0nH8Wo6dPYqYrsYzn9JeAKbSN6j/iDMtJRXdEczwpMoz2m
dPvj+NT/fXSpiwmAr2hRhNaQLEfijDN6ibv0xOpdWit1VTmW34s4LRXG4KCJ2OfIV2xg1T6jfRKC
SpZFSEBQ0sNxo7TJfbAD4QW8XGKyIJ9xGVi4CY5H9ZB1qzdRe4+1xO2PziVDz2d5iZnetbiQK9lr
B7Ub+3LwWQtpfHoJN8QIc04+7h5//m9aaBDFIwOFrJ/lTm/3Ua/uz9YHBogV0T43qjYjGHXFNrm+
3AoVhz9FZFDSeZ45IW9mS7jvxrn3KwefRx0TSWNs91N1PZlFAJ/XJJn8xg3ff3HXLaE4YJHkw2wk
IchgdR58LJt3KxTFYz41U/ateErqrktraRFq522nWeopiK1o+49BUiAnDjTXJyuNZ8U8YTYeo/ev
COSlM7qDN7w0ZuaABmeGhOjS5Vr1PifVrQvtsGvM43RUyL0E5a555U6sCY+XgD+K0nk+sSysRldS
fveERa0M9sCcM+XDjmYvG0C2Efno+B+ALucjsGzEGsR3Nt3ldbvZr4tCl6fpmv63n4OxBLpFF+Xu
UM6IEaILScx2trG2ArHzjgGmj8fLNCYP9tN9cnBKnLOD3gNRU22+cKtC+IzYrRh4vW62J5HYtaOH
5Js3WjzRczN8QHobxJ0Stqf1uo0NZlQgYG6oz+qQ6r3nonbCC6jCrGZwCQrtZCHPcfDcNDDrhEKI
gCm5lQYmnav3mTEv2zbVgL8IUTn4NICIHsgRn7ip/0KwPBAQwK+V7Yp8TVvVjKKB7KrJLuZfGrt1
zV5HH7R/XTkS/Xsi+nWXpVEWlf9B+Kv2mbr6jokFvEoy0T4ENYWJIKMLZIf6qoSqIq61YFmYxmt7
w/wWaKWRDyqkdJXQQjklEE+Sbw121hdKobTbA0yO2rhf3iH3tSBRVi6nzXIAFtZAHuWlEQAJMpQw
TMoCB6Feqi7WTivyt/hy2evMZZqTa/DFKNGL8MoOoHh9oqKLmG2uqsTaDqoi1Ir6ZkSdyHDa7gQk
AIkvjTYk5vdrNuJcqs1823VcPZSX4WZAAME9usn4SpYd+asdYeOig1nytQmSvO7c3Z5UzORWGJMX
tFr6t1MOkBYvytOn+2fOq7RgmcFgBZSLr4N/feNvZW1rKQs7X4AmDPIrGeubRZ8fre4cuHg2wvKI
MX1Q11lbulb0iNqZPL9KJ8bysvSbOWCxH9zlDuiMvUUEGciQl4Ghswgv2v/9e9IH3ePc2z12QW/J
p0nIFO7/4qIWbCYhY+dKTrENwMy/fze2Xp0jcA4/uMSDHWVakiafNh4XeZzg4au4YJlYyfXDXL9S
rWNqB/TABVDyQ3GPK2xFiTpYQH/PsPxowvs0cpHEZZ9dhBAdgE81esIZqeDcor5gBSchXt7s4xDk
kXjshdIKXRNQbO4y7KMeZmJ4REbuFq2z88bJTX7iCzkg4KUP+ZvZh68bqJt27JrZEQb5axahVb4f
3oexff36CoEWUW9Z4KEgOlaa3/fZCvEMvc3kLplZP9x+TnKnkx5CsdZhidLo9gh9gPdRKIIeYMGp
kcOOP1Zg3mG5ZPafkjkjsW3NTbqvXjIXpx9L/XY1DlRy+CND7tkS0SQRAUcs7e8sEl5F28gc4uct
c5wlGYMAnQVWNwR2icR0fXeRRGvKmhP0qZA+yv38yqsWGbCpOM5un8BwAe1JaXCAcwmEPcRy9EvD
WRe+NEglrb14+xBZpXCUOLHRpDcjqpoDYZ8/MM/oO0i/3FVTOLMKDm4AFjGRafswU/ARZDbrcS+b
kyuFZE2swnzyUGBuKZ6e9O60GWVlSO2X5Ywuh+QCKDZXH21SRfRI5A1bRanbzsmI6RolBDWkodJp
2lUthmkY9lKp2u+XS3uhhHKWteM5AeDxIHuV5Lu/gsoygVR+JNZShJ0iIOhXroxl3gst4Ik4RhMa
cLVbI7FslTyItAWmXHGZF0dDSmjuBuqlH7xKu1F816fMjCN4Ul9GZRPynr0zxQX6mkSPP1mYWcGU
T6/CliqbgjPqfjpipH6KL5Tr4VXZLFJjnsijv1gxK4jOm2t50exzOBG31C/LxQoGA2rXFSa7+EAZ
Q6HF9kDtkbRMajvBYvLbwc4m5ZJVjXrjhUdsK/Y0SKzD1ZrMC+OeVyQSpipYjPYYH5rohkNJ//28
PAAxUwpRGLifPV7F4GqYE0mhTXNT0AYAVOIP4NfRm6P6qN4ORDAT4A9SucfYUKP1IZ2ZeAR8t0Im
G08ipA4sVOybMSoSjiMsywGDTLNNLON6wixNRFm1V/U07D5qNmFTMuwcyaudcJgSy7m/EoYkekpv
ugeuVwc+4bI8wDmH3+F+7Ax1IVha0H43/84R1c24I1q+vlHkdO51gjcNk58+OnuLRqtAPkiCBM/6
IXgVGRdt134H3Lwt8GAhl8NDP8kaCQwyp/YYXyKGnNFUfqCmlHOPz0ttdnN7yh+EP5rqDcoq7wbK
im86/Lcf6Tmqy28BAxuZfzARDcGXLVvGOB11EcO4gBhWE+76Ik6H//ygejX7Sy1YTe8yIoGuxBBL
hLI2w7gj8QjR4ZW7EvWErRexgdR+3FSniCDJWfYiVxJdSF1MD3/dL95MOGApL71ZZ3hqmGFQMwyA
4Na+mFnHdcehYYJmdF/AhXUeelQfJw4VCnzEEIBh4nFR3PO4W09lUjLB6QhCLgqfL7293eqWI3e6
nwx87vaHvu7GtrvIZmdXvJ2Ss/dYWytiNIjrnNNUiOmqglUTdsNaaNd/e+I+dSFp2XP3Q9mBZtGO
T0Glcss4wDLsBPPi8wSyxuJoVl1RXg3PnAEc9/2ymdj6Qr8bVLzmQoLj5UyDP1udEJ6KAwNKk42q
07s21LLRq6VkxAglg6Oh93dw/KBC2Iy1EB/YTyLwmKn9X5s5NZD4JCklJ3pwGbD6Bk1W2nyZLO6F
ov6BNb21TYVPH92aktiiDdCRXiR5GdTG3OC6iXLZbmtiHr92zCiRH4dfB4U3PYPGNwhJef5yKXo+
fhHI/hi1uk7hAe+WVTHL51FzDmQx1pwl194l31ZBqhRDSwwWft96LOzCcBIw12TNcPG8/H/bYKA/
SCcTqUAWl3xQT5wBrs49P08nj48ddLy449SdONChzyRbp2236UsB+v2jGlzOkN0yeVlfLRk0hrbw
uNTjWh6QmmZ7YA7mTLWfKQiCVqb1j6OaklXhQCq7Wm98enaVRTd/tXOCLLL9iLPMeL2N6M9hgJzs
kbrWGUpGDZcD139K8NASD9MEO7rI6jwPBnRYTM9dqgGYYTMs6Y4SXXAs7DsdfJGSbVzHfjLRK2KC
OqOgGLWDOdmpj/WWneBaCFcha/JLTrK7uBbF19LOoHXpAXtm/TdcKhn6P2RP+OvK1GlEEWxPoJOH
++ga2Ogg2vKuzyWrIacJ5jqb+ACO5mQldNueeGla1JGt2RH3f9Yo17c91FFp0wEjHYUtM2Gz69fb
opS7INPi917Q3gDq5ws+NUNhVhKfvsUiH0Dd1wEYaXAWBA6SGHtp+aMuPo4TBuLjqoGiieY6CZLA
nLPG0A2ifQX6fom3DaSAFVUE+Wmm3du9O46v31rH4ufJk9mC6LPiCFCxyK7seYYrNcUqWzhzMwsm
Mko5rhJq01PzvTg/d1jExnRJPWyKwKSZiCjZZWAvUObqn/2uslcwOX+RLxl4uAjJbdfLfHHy9auY
mfP2MVIfTH3Nhpxizof6L3Yce63Fa4jBsHUYRrQy2rvabE7SkQDoZnw55U0LAh2d31SKxtBN6gZd
/CycBk2L8/oTuqlUxGC9GmflCsWRMraMkFODo+D4I6QuiWtpS4+mc5aKYYLlrLK99zT3vFV6MO2a
aEgfRmmRXLU33fmFYRcrlJrFr3x3oY5ZVTWJcCEgrSXnsvp12uaUMxLVoVqOhrvMIObPSPD8K2AG
APZaveQETPdkgBJeN3MAANn+kKmOiKsWf2Pppp4RkAuaz2f8nVfvaZ+NrRIysJRyGfC1I25BCg+D
JIzdv4SdVNk3QqGs7qhnlXN4IM+tN//hTVij0BiR0AlOO2iVJA0u1OLDNMUi1W+rZGBjBWSGTzn8
3zRDapdVZP48u9RZ9nrWHJAqG+x3//fR7JqFhrPsEYBgRfNBnf10UOf4NZaHCnJnftFw65jX4Aqf
xY/b4Btpt4PbscZr5EvMz8o5INVoLWgeZjlvJbxT0OlEnCv7CZX6EX9YLbfoGfAkjqR+40qukIsB
lpF56MOOJFhm9goGEJvL9Lt0ccOCYUZytZWfZEzfr5SDunVthFIqvqtce9JMKoTJ8l+1kmX2D4tp
6PwYtgGJJ9VRWjBh9UrDa3Cfcej2rLLNSDYwZAOJTV2lf/rcPyPzrgTZijUpRaxiEXo+F0M/LtYA
kDgJCCr99j8K6/C7k9m0mkpuJKFpy1f2reHIHD874FKw1608PTNS08DR5LtIhk6hs8DFpxYxBHaV
MqC3Zht/VVbSZXG9g8+bYRB39qXBsidh+mtCknF4UeiebaNrpbgDxmgsjBb+zO9PWJjBo2YRFpo9
D483l/jOUuouECs2fIeSP38JOPiKLr294ntIxQsu1fEWGqRxDRqLUNTdFVUsv5MPDb6nfBhPjpo/
V7Dy6AXMT30VY3K6mBuRb5KPQU5Qlit+M9Hn/blz14dSPCZfItXvK5EvzeZUsY3TVr3LJBGZzCd8
fAnhz2Mr6de1N1veYqT2SLq2c6cTojlVuN/cx7kWO5VUDUGU8i5m5hiMAcyIhGfYovHg0HqpBGMg
AUlPw1+xHvr/4e+QYLyqZ4QTKpTZ9A8AUlDMDr7nXLyCh22T7frGFPV2/dR+CJMiuHQxY7ufE0A2
NKubSbk8pt9hpeP9c1PEBEHWyqoExczCdL1TKGh9bBijzbJQnph6vglNbYWAJrXHcSaxicYu8C9R
8sjds/Ugx8f0fptubGpQGU9b1kR4vHygklKO4KYuO+2CcF1TmM6clrsIfnCarFXtQBAGti9Ix2vb
ryivEIlSFL46nYovTKrPzydRjpyAS+xe+is8Rk7OXZDdxrQ+nY/EjHZD8d0iD3AUSHSmNSmIMKZz
eHoDE8fUbc9HMUcriNYd/W4BMGAsxKqIEaPvpWfktYTg7OKP6ihCDBRirZIeB0sZmoJA4DirDN+F
pigCRus7kj6l4UEDRqU8m9qtHpiPWD174WDM2HgzSULnplGaXwC795pUj6Q7hSKOOGiUq07Tg4DU
dZqHIz+V3uGW40FxZaDrZ3oWsH8quuhM/lxVhihO8ayr+YZP0ImfN6RUIFysDBn2gKaqu2V+GYMc
Vvop6FSZGgOSSUyzYLNPbiJ9yvToyS70PlOE6HqewT6YOCtjaXq9JLzaKwg78ZAAmwGslwNCXN0K
T3oTAa5uys8AGKoCOpqinfGZLe/EofpIZZZIvL+OATEWzj7IKmofwLBCq83LDFIWbgzqe2hdLjCS
bTBEIbNn7BY00e6Jsxu7NIhrRBrwHatfcTUE9yRC/LFEG43aSd+z94dnbOEncEwYys/gEw5QIdjh
ctVAsrnwYF+MDc7ujJeAZ4X0PZPPfuawqWkiGImHKQQjjNgSNzVX1bwd7LgWKB05sOyJCQ/jl4vr
Z/aMWzDRL9zdGMxchGcQzHC6yhkde5yditvabTTM/61FAme4iJwmQY05TRMG406V+HuTZXxaKuth
JnLGFaJ1dMm+kccZqHG7wpushp/AGLgX+DCvrhDH/W3St6JTEXw04QThfk6Bqr+8Ri7ynmIoovHh
lmL6JAJ9nmXMjcPl18FomTebfcAuGeujlyuDZkSUjbz2pO1/yoIDBZWTZCrDtBt4Xd0Gq+OpwJtq
F2pNdpkO/Lt+DtRaoQyz2hmnCjiL54M6my3dH6d7KroFFWQFiMSWLKxUQ23tbJYyiOT5F5sgnDls
H+EMG+CC0x1QpmUog9iKovUcch/0HB9Q0I3vGXM3slfBu0qOhbNejxQYE69u0QzLUlVP5WkZhYS0
U7Ojhy1wGrWDykKOa7gDDZu2NRbmARDKNkpGhPTvvBi+9OJjp/NghfvFgBfInhmzp7tEz8k54Yq5
2PdlT8y/pGNOKMeTJeR6/XrnZMIEhtf7EHQGHeqhQccPy48fvUe7j7NeSN2aCCxGcdBqPqTpjOYr
hSoERW6lM6ZKv9p/wz4NGpd7ODPnqbLSR8rBKtOo1FiY4nBhPsGRyGWNN9HhWyWvtERbbic6PCfy
mrFYPocTunp1qv2CrN9iHjYMKJ9Eo9pgwkDZqtVnV8PZw8K2NYUDnVksMjS52kuys/U+Jz4ZsDPz
wruEZbcKAWIAv0eRZH+hTt8pRhR8/OcsD6ZAQxzjBt2Ca/r/NrnxjsV3XzuwMvceekGnnRRZ2oHx
sDX5rG2x8rCaWCXZ706g5sj6GMrFADH7oq8no3I4L7cOjzm3jSNUoNzorInX8GjoOjqlHPJoKa0d
NXFCUnUo8yTTnNSyNaLRLdB+41tuDsO3SQ7ho7if3zwAmJOoEAWBx5ZnNbj6bzgDtkf+NKI0mdtl
yiQzMabbQLkwry7P17H8feLWQURJt+wH07XfZZxmRpqutdpemnxa1o4eJufJIbNzY/AHel3LlSRx
e4vACo6AvGBSt9g93hxZC+AetMs/qoycZZfAnjZnam9t86qFQpHvcwcHeBTAqSlUAqnRo6platEI
1XzLap7AXwUd+gqA6azkKoHxrAwPrxvZPL+IhZfa+WuE0VlQ4JX1TMkdqIIrQdk0xSMsJIwbhtZN
S4pQ6QLcUBka7cflWDsa/SBqC1gtmFGI6yAGrazBzmm/CO4zhTS3X8VwrbcD4wCkHCPzspE4Fx47
Yix2hrktteT5XWoNpCQrKrGBQg+ga3Uj7CSvsOfHrSh0lKZJCpw6rvl84JeCTMSTvpYRnTED6cEH
uQ6Zf12ziuXmKH6sdCx5verpYtRzrnNd+33u+DwudYbbLsGKphL8uWvdf/A4VqzMRf2oxe0CQBl+
kjIblRCALSfWPuHPOhtZywpvHVKcRqgS0tR0VcboE/B1eCfFaNQHhVV7MkOpxrw3uowKvLfl3LSD
UATSukgLk/v1HH30T75BztGpuj/Dgk4GHF9Osezztrkr+0g0b4spUvnpIjiSInbenjP1eElmHjCc
YokPN38H4E3gctBoNqZksma5YrmNedKEbhAAzd1aPdwid0bzZX17yxY2c25yQGd9zSZX9CxlYb5J
h7i0Bnhr3F6HJuBG2VNfUCWMU4UcTxnX7BrDV0VarovS9Gqg4xjhA+fLujVhPC6JffO2N3/nmsE1
BPeGkOwyr5RJfsJavIp6SMnV8Mr18+NaAc8vQoBk+viPb/CgdFnqfbwnRU1KvDEamsaIGtffnnYg
8DT6CiknfRRiCxhLLaDMpXci3llw8aAVI8CO/FXUMX+oR2DUpQsMNote/PSpyProyajYgusB/vnN
UAgV0zeYDufAWBe5QkYSF0BBIyJmf7GdxJ/+7mwGqcRx62hYqUx/6VR4DxUz111ZoArA4Iu2xtFm
UgL4XUtUUplmcYCOpgEHvIFcZpCXNusL9SvdCyel6sSW0Rj07/+CL8D0m42Z9Gy9MaWV4f9jdDbc
T889PqK6YiFkYhzhcFcNPoLWm7SdyInhib1oSEDz6Nr3Rg43RK92xzA+bbCMWz6F/xaW5nHL35iw
3H4pmSsqhr2q+BWLPMINh90fvhhYSiXxYpo0T0LgHfehM/xaLM9LFUJFpL85KUWDAe9+tcYMkaBC
7Lei3P7K1giKBiYB2Wcybj5qhoW/YlIWTJLt0HmSMHaQmjUH99k116t5YGHCJ0QHz3BgBW8jBLaz
1tuVU4dMnQjPjP4U4Jqdb9trAcSmeCdJbBEHIdC6xNk9uLdtf2d7pdSiyuzQxUML5IPS/EQr+DrN
xJtga7aPUNHzyrMrSVrtyRdq2t1zuGnhTHdvqJN/S9R8JoHgfCNtPA8YxN7rEbsawz5xQSnj2urW
0DM5/vNGlbf1e5iVFzJi7Z5DWefNaCEUwMY7I0uN3nNRdi7yaFpTUD+Zg6j+NDNzcIH0keHSIsDP
MmdoDHaChdcVlDbIvbiB4jcnRYPeBRCg5ZQnetLhk2jIt9D3OFhWUNoFsg7HlGS4LeS09gf0NvoD
PrrFUkT4ene3WoqUTrV56HlezxPozciQEDfgQiVUcliFI2J2Tv/CeBBKkLk5f4OxT+UBlKT+eYrE
XfwfT4ItkzOhTE/5HFNNyGmzetXQPSVCvaeU29WwbB9H+Oom8MQ4kBbpCDbv476yOX9kv7W12BDT
AxDCQbmqjy4PsQpQ4KLaDqflTtVm8XMnksmAJ5xNugd3Rb7ke0XetcsQmK0YjM1vwiqeeeQ56IRS
MdXA0p5a9TViwZMsDBz0zqAYj4UbyWmqHrACODwJ/ZBYorUht2n9gDxZQaTPwkJKtzqXfgV42tHv
5B2UUiNF1xOg8YO+DROVDyUuC/gj9loVh7m0UMOSDnD3QbADJRgsDuzVrAcaqKB1IGPbWRh7CPZm
rwGGyiXwBfr2OIGZpVE56wicAeu8LHowAe2gfm54UqdKYHorPN3ltOogmjiKs8LVRLmPS7Naag8x
2O+YnTiswmSoBT0TNjfaKPmZYhfJxRT80W1MCYd0ziKENZT3PfphmjzQHJDygr+NMWE8e2kCxNxx
yYJKjp4MlJcy2t+6c/3Ybvs9e1p4WYC3AgL4q+CsYo77cwQeIi4u5bV+fPxBafB/nHxh0nDYEHBJ
UYTuAqlcYyc4JBNV2lynb74aU+5n6JyXAANLlm9J8s8UPmSneSOxG64psKJ4njYFRi2ny38TZAS3
6Ulqt9RaLZ6mSyFZSB7Q1RUdsHmOQJAOECYWS67x9qnArwGPQpTCPMQF4bDmqpG94LdmeNle2ntA
3XqgyxqhuDK2L+/pAue+y5w6wnOcklobH5Pq81+79vYbO9+qdPipisBO80S/eo6VjuNbzU/KkYUl
DUY86EwE4uJ6mSWFNMptjoT8/64wZUZxVvNpNqzQvfZGyZU8KwFw5ITX3k/DoC6HMb8c3EozHxbl
l98u+vPiX5NHUcpw1Z3qZQiosDzytSr/lbiNGOjgGmt67D9gwJXM6GdbfglH4yvc/MHUJ//GCtcM
WYfwRA9EHGN963v8C3JZO/BQqKHpskEMMwkPAN/bwkjb6oF9QdlogWFnkZHJPmgLNIgo2K6S/lNq
kQQxieUmKed34m5BQPvu/nit+9CfRCOK6CgcGEbRXELHfgXIxWFMY0krd1rzFRwKtbHrmxabj/FW
XLXDmjxpp03fP13+h5GK7nw6gdNsPSMQagp/PgIKzAZYy0YcYx60MWszGBFRjeTqhgiTCw7HjlQ+
YmO54cOM4MPjmSUOzVBGXRptrgNGX7FHR+/0SeVUzZ/IBM8nce60xS2+sWlDoo1YvoExH2A2ZOxm
Opcw0teAmgylF6T7EEerHc0qL01/wFVk/6/a3AqCXu23vh7o0gH/2cMMrWyRtVyai8DsWWnbnkc5
U+7Sz3NKi9qA6SVcc2QNvQF07uuQYmTZNqFg4SbaWp+k94jYkaAtCeS0QvraEWtJmQYVz1v1X63V
o8J/5dju8orapR5og09hM4V1OZpcoubYBDgnciuk1u9N2TypvV9nkBUu/Jv70omXXBwiNmu0YTVX
dWNEcsna4mFF4K6gezeB0DG7PZ8C+WWzyTj4BAel1QysfaAF4cXwbW4qSJxs0+DX410VDH6WBljq
uFR1NnMDt/Z+AXHHynZxvSK6dR9GUPKhug8DEZ6BNvkKgiV62YprAlooyQG1anrZNQlg/kbpcmYt
prMc67GCn8ETV+zRoQLqJazlQ+TtZRHuE5YWZ5kvcHYQrDdP1ZyFTHS3PbEdfnsSJwJ21lil4bYS
h7jLNK1CztSHWgvFW9v/fQ0NVf/kf9KcrQznvqaDHdMPnghwzqaTcIMc71d+Or5YH7r1pj6d10LX
Qg41RETzIYvpMO8l/JkQG2K9SwmGnfG13IVulY+D0+geD7sTrMugZSMcO6UBYXkAMv41ZXZWhL5Z
E9dRQUPc+vJCkuzRGWVrxpEk7wSCiPKGdpzQ4CC1jKjwFCYjPBxDktYraxsdD58DHtA0fNzgVOdR
mVxSFQhEpYhYQRqO1E4gjyvuarqlhFGzzdgq+TaLQUzRu0RIHlxS9A3z2IiPLttMNbhOVqnIAZog
CEnCEIUuQhkceeeMYRlLhuf/QCdyGrMmXfYjqMVjPeMwfc5wDZe5TOMCrr/y/0AKJbax6m0jNOrZ
haPAGfDZsKXVrJ+GhLGd4tqZ99vIBnSSdkqz+xsA+90gqfnJ5omuCyhjVs4OT7NRn6QXSP1vD/uO
RGpYJuLh7gLYBKNPo9nQylw2nmfImt+Mu6XLZGt1GIaA9SwQlIlVYNV1FdiChOSw6nTzkCIx+yZo
VMCxjrpLAaK1/N9Sm/tyorbpODdETXt0voLGHIQ+jCLQu7ZsU1wBV2Mv0+y+wgQnkzytplrk2Byt
J1FK2SeJnVic+wNFcBiA5Lns5uOH8Lz/gD6BD4brvftFugZptWC3EhbcMMq8Uc4kzaNgq1bDDmmI
v4IDGiuM+eZv8ZVkN6xwJrfAkU1JwtUOQ2nIbpKpbvVonJcyN6o2BGbKD4bNP5iCrcFcF1gQM1RV
LC8RklkU6GWGYkpHHSTBfaN5RgifqADA7kIMf+UtYwPJbutUg5joIrbCOGHn1o/PS6oDAISLdDh9
iq1ypBG4xCTwygijWpBmB4mpf+1Sm7BdiOC6KuzwwnQqXpgFzGIpx3nyvVchDNYoGnma2v5sxblz
3toXBu2/ArMc4x0IjKGtgSffts+RyofstdoFZ76Qfte1bP8XrG4Kkbp5Mng+qor0+aQIR+dqRYWc
NVRk/LvyH2dPoevp1OzFj9JjW1U4+Lv+ADplxi5i4AnOB+fCTHl+mSQLzYlBQZ268nP/goCJdBAM
5Ma3FIEmbig+rmbVio6wFStqAUBKR2a5LEb5NA0thGwqseMt+qnsEtRoZjMQWMGjFjPh5bn+pIMN
xO/jyietbuS+DF3BmldqPHl2PTvZbUc0ztVFU5Cjl9W8UEY4oWPj64oAQ7yJwc5wuiAKx6is7efA
hnpPPIN4ykxe5EaaU4YICrrAOP7Fpv3DP0B/4xnhXUmxivjbtIv9Z0Y50/9sNEvMbhE1aZpbe3W3
d6iip/QNsFlfMuZQGOM8TFNB6SMf51CDOslhiPlfcDVsTxgmFWnD1tg4jwC2/itAF740VDCLmTqb
ji5TLXVon1l66nETAq5cxvg2Wpb3W3eIXSl+kcbjm6oUV7KhQwyLLK/ALjw9F5HSa1+t2LQIT76b
9yaXJxxKmnKD65ws4Eus8kQiQUmWgnDIeYPfndau3A3S1ADd+lwOZP4bxq6ylL8EnpyWU+yM8u0y
mhhhy6qsmmzljJ1EJm33NR0UuZid5Q+sxRt2u5BNkdCgdiLU7rGTOMwGMYtO6rtUnIYagG90PYBp
9slI2Jw+NYZBhESq9f8gC5q7uB1BY+hbaZJZCt1dw8afnF1DRjeRudM+e1az41sMFDgPHbDR/tdO
V09FZ7x9IvOq8qttMUS63fkb7fRr4J86EqB5nuQ4qrD6y6xoe/smTQvsWWtjXW/A+q2g4Kn6Uouf
nu6Uqr08Em+iGxU2X2O/unediWVZt/rUuwlWJjhAneuU/LMeFAMGrWwjru+pAudhqsBMlQafMObL
6dbRteaaV+9bMd03HLpEHAD/e8wnRY9fOyxCUqGQK0hCuKNuZD0Fdei6TqgTvhFS+oKfHdbUxIbV
ALvnJNXi8PaBy94hjuUVn+VBtfOK3nBE083L8uLPbDdARo77cg2m/SH8B0XBrvsDoH9shbOGS24T
UOiOq5Rtw4gX075sB4kGtUzKs9z/kW7+esEcOzd+BWfHGTPcpoaz01lZPs7yAXaYFF12u4pDEb8g
ZlLwkKsg7f9SdUE4xkw81q2DLD6P81By7bLJSE4orUXAlQlaUwmd5EiQBONe7QC928IIOi9ZfkZk
KLLXDL4LWXzxUUpJFS4A2FjU9bBqRPiTamIRfrYmmuucMtsFdoou/oQfJOY+Eh3uIdknlGcsTJ/D
ysvo8qRAUPSrTbJCztwPB2qa5mxwbv67CrbHuMwE3bTYPZA5macDThy49s1AU9wNdGXQtpbLZ5xm
BxQ6Bm+qPvSiwrw+kvuwbznw64fKah8Mw04JrvmDFTJy3X7oB5acm7SR6Lkm5CoRRz31n6xTe3Uw
xDo1aoO418Y8a/8X11hvoZmxgDraWYcJXaUz9pj2Xs+VGzrolbxQzp5m5FojxPKw6ikMYoS/bqiT
7YwTo+C1dRsmnASHpazz4kqKeZFbgvq6TcUGYskPOFwmgvfOaQpFTbF34HUASlb6XB3b4ZqMWlQN
saoq2ViZrgUt/0XKTvUD0/R1GhmQsMrf2sl4pC4nU7uvYlXW0nGZnQeiPe+8dfrURJvxWjNRVWYu
KY24u+q6Ho9qEc3DfGQ+loWuOxWyYAYWeknlI5FukmQUOL9x4y3/Uz0IrE6kdvzJqNrbhYYBSzCD
lP03tDA5QfP/ohyDNVVYU65oO5VdINT5BcPkUhPB6+ca0ETjJXuTzkPgDIH8x9l4V0JFp//DCKcc
8rHrqcoPAjJ7zq9v50awFO63Un+UukPZyvjuYvOG9msO9tE9WXKstGLA4W2synzrexcb3NnUumqy
B6RCecVIWwd+qLAuRPUEgKyutCA1ay6rsVOS9b2tcCdQWlNf2mZv7asuO2XT6VwUjR+0mMVNDyFG
tgmiGKqrCKMECZGTXTVJtAEjZbS/rfegfgJuBkP36lrpzoIpT3orU1RwvLdxWsw1U+ioe13d4PKf
V9rQ+eQuNVQIJl/IG7IoSpK4MUEKfpJ2N542uw9yzPOE219ChmW0AJtjnQUoJeVUgKP6RHNXyvMG
eLOO4/y/UZdU2EFuKzViS8auQHenmDd2IWi6jUZKJXRweiCwZqjSiD1+BuTzd8EyfPlWV/HNnTzl
wc1mEHR/D+j3XTkP7aVFPv0LpHW/J8yB1OOphqGe91cumvN0g0H/q0O/IGPPGkZ58mgpyO15UNZb
qJS+D6Kk4YDwdlUA8o/+z9kbJZ1BBckHaCwGDnjW6+PGZ7aewi+4NoibrdIS1haTH0/oflwZwLq+
raJ+p0hKeM4qnV3vxFYAiEwEZ1FpLGUOGJmfmf5sxSbi7gBlcQTdDE+E2QlIvcXKI9HE08VKkljq
F2upyFL8XcMWjIVNoyXrmnwPpwuyxbF5446XmR/lmm/gwyOArLqjnaAe4N62Xk+HHoAPbGY9779K
rsbsazeKqGhhg0hjlF6UZH2hGtfFVTEVXLcy/IClC89B28nUKbdFPo/wLbHBUow2ZG+I+aTQROlq
HZ5gEzQl++ti5CvkCwEK0KR9I00Y5naBK8z8o508cqSkqmWOmNrrfke2LbX9iUIWq6Cu/Mh5h0qS
CBhCB7v1hJ6fwiuATHZ7S8N43ucuZa9AKyYoH436Vy8qrycExD9Wdy0alMLPtTIwvvpxh8xDFUPB
qyWMUJOaUCr75fySqqeB4aa/7Hzkflry0VfH+VPH4m6c8aGkZGGw8hQw8dlr8bnWL3wi6kIWsJ7f
RPTPZQCBXTVXb/b55jKDSTjPRoErVkW27iN976jJGUPBCLDO3+ysyAeC4GoH0CVgORGGaPMxO/J6
CF0pWzfMaJ/01+UdqU4uxqpN4DbQVjdCKZbiYQPmAukbxcXB7MNGJZt4jAcWOQlkypyoNZB+wtwA
PdHseDbrzPYHiAzC5fh+DDivytCqNIBKDZBSHnhy0sh5pcFU6QIv8RMmIZVwR6qA2Ie+qjUP+ZzV
yrV3kvUC3BhKm+hAShkMXEFmoTrkZmvKGL54Abd+jX9/3gtQ3/UwtCHJ17llkhMrXFnL3PoUau6+
iw7lbUVvBVrYv2TFRoOj38ctkiVYXgc7GbNykHpTUYc6rwWJoUixfFYL0s4l6fsdc7u2mntK38+u
CgWszQl8YXUMH6141qwaE3dsYb9PN7IW4rJJD3IYUOiYW5pqPn4X6meTlu0Fs8ygn9RheeMer/fw
RlJKucWrvsU6y3gPHvALl0sYhqfVnnLmqtgeY+x18k+xqOAdm4e7Pu4tw7uoZD9gxvbTZy7S9LaP
sF0H6l4M52isHRVLbaOODT+aUmHy2hhpDcHY7plNxOthgxVyFUvJoOQ+M3aqIttzK9laQqKzbK1M
yG68IIe2McXPqDk8Q1BBAsobE83oiOis2RVQ7pvX5TYPwh7z4omkBTN+DJVuyjS9a61glXmd3MNk
552hGGCor6BfwT09J/h0mCAWbJPB7zvtq+Ata9pdw9CZsD32JMBX9sYAegiT5AjiqOLyj7tQ8pU7
fkn8Bb5nzLJeBU/xZkSjJU89JT/TbKWoEC9XROE5Rbb1iGpHuujG6IB+qe+pGT8E70Abh/p/oZ/Z
lGZFEJUSJb8KhOY3BRHej1HZOy9t8eTVozKzhSyHgHnuUFFyd58dPjs8vxiAKdwXGeVg/BJxZnur
PnZZUxEMUf2RZxU0XVJNajLMG+81YZBAztgHcBszIJjL+eUYaE55+7vZQdhSULAfCsAgV+To1OEy
Sw2emE0Vg9xx4MPvM5ZFidmwVVSjLT5pnE5F6x2y6ngz8ejDuPUhlloCUKhVVowGyCl/vazU0CWs
mI+LrFQ9EcNe5WY2bk2rEkk0TmFT1/FnvO4CJphMmknqSeO4XumgtCBqzGBvXl+ZP7CBd/ieOPw2
XwMybqDNQpIhUlz0teqmKPzuFCHGqBcQE+6yhStRDOPsp3VKz2dQJV6NpYpS93jOM13Zdj3NSwS2
OhMsk6gpMfTeSxlSnPc9EQr5RN0Fi5MPTls+KvRw5KPb4YmxOZlCvWWHXblJl2QGeiI11z0mpoeN
WevjWo/GNgIXmBCxwbd8v78fD5/gIOjVopcRvUf4w6jaryYurt92VvsDa4zZYLr14eThU+7F7a1N
bhz7NwgzKhw2BcKDvW6NM0TEoJ2pjOMZMgzK9xkFIxFbdsvxCSi5ryphLWVpPFC2bAuYuy3d6MOk
oUKEWF4JLIvqj//N6JfEjgDZtq9lGd9p33Y+8Zu4VV+tXm2dx+3CBTtjqWuN0EGQGOCUaOtkphkG
o/PcSCZhNDmIhoudwjIpFAdS6DSHHpDRsc+hTHKbfi0CXTSsYOutX45zU2nATLCEsX1O5KvzGF2U
7dosAu/kFPXPc4suNvAetirV61a+87YA2LjYYDtwCOYyZj+3mw8Xu5C1714XqJNylek9wRoeQH7L
B3vg9QCc9+gfxtli3Bp828mhrLmB/8ych9dUTVaYa63P8oe1BQIoP1/dmXZVu9xnwcVJMjFPjtMx
7UiX6K1dGxvljrSdcWFpP9zpgQZnLGz+E0Q8CGSeguUDoTzDOklr+e+EJ/nkdS3AZU9G6CFs88WV
3PgdhkIuRPx4KoO/KL/YXR9Gp6jvlfoXnMDKuagACw+9lmNCRGXBvQSaZkoQGQ9jGW81Bcbfxcek
iSsb7iXsX4JBGoPLJhEhbzuYhGbiAaUYffOy79Xg1oEL8I9T54KCf1drFT0fZDX0Y5Ji0ac4PytL
3SnZXOZGvjc34tm6It0iP7L1m58Kd5eI5f9PQsaxEef0NbzeODP7t34ZS8hgBMEKuy3xeCOADHtk
jFaGHDlh625iPdcL/pj/lND+TA5A5+KVgbWcT6116lK9FYpjbZ/DA4q4vAe9Sr1bwklWf1ebk0PG
eviAUGdecll1xIsXoncpC91rHhTAD+Li7YJ3Dixd/J5T9XRvNA0gM49uDQC+ShsCCo0NLdKsLPFj
si6QGtfzfVArk9BhLQ076Hx9hRxzo7j8M9G8MqV3GgLsdSHBD00pRrIyeE6a9H2rWGCT3zTMhmwr
va9qPFsou8iUZ5Qp/E4pVpnl9kIQUpW8E9iZjRjfanNA2Puv7UN9J/vXi3mIPOGx2Mgz45XimYr8
YD1SPOCm9g//KP5B3xYDf22rOWGXNkfFDk9n2zM9DCbS+lUWEqBB+YmVEKODezTDDcOssPIiVFN5
OnNbnMzNIkQvoYENc7ewWbuaDvySlb24WbFPF0hYfhQ+KUNzsopLKD3FPU99PGShpcX5fit3fCMS
8MNwQ3+NaG5uG4H+R29dN7xwNKgFaQKhNxKQtgvVLJKd56luT8Ezs2zIYBqTjhZ7CU4SCWgYqhaA
JQdqYbw9UZWRSSUqnwbIUV8DPn9Lo3359VbSPS45LYl4piViaSxVui6S6GScnoZyX+GcMqoihRLb
NaQ65GWwTu73ouYdL8hJYhUbJTui1Kxx6xHaONig/b1eKy5mF8bUPb3xzhUDvu4cbHCnpL0Ddu5N
zmRi2YBVVh2lLlbOc74gC+L9ebV9CdEP3vqq8Vfut75LjOk5i7LaAqTNF5SWj96sXk/NESk3mRl+
ubV/gHbc+3AOCb2wNMPt9hxyIYC2z79whXrW09vEKHgjgGs1BPpU5tiajlXqIZRVSB20875Risri
+w5mkjwVYQAQGNzQtO21EuP1JjZ7uwcLtnJmRqR8mS39HY+4wMBYJYYxAvRzKi9Kp8kekH4sBQik
0P5zjLowIiQSwRvvWj/VOy0B4uLw2NjStz07E7/eV/fWREey14j95XlLVwHGwFwHxdk13Cw/W09j
SHNXQr6ZGH/MVZDQz771CZA13Zpty1vovpSnI1WyZ81iDQag3HDcQ73yPI8gzLyqHlX5ohmtr8P+
5yVZdsKxciAa5l17TGLvh5ZOBPJkJIBNWDslZLhSVy3lY8onPLcyWnC8BfXoam0IlpQSvXiF4HVQ
/E5M7ACslKfZZStJvmj+fcW0HUkqRrfg/sdSiEEcsGhM21eNkjeKGTeA053E/6oiUB6mfarYQ5n0
GDhn3CvEXqAeGXSMcxf8WzjoCYAANtAjWXJmIS9rYr2/ZBYfHKwGcT5qI1ZINu5Q+XVsal+Vo4Fj
mzA2FP3TGE33mWsvj9eIw7Jq9H58wnEt92+GNwub/mwKiryOm4oISSSRxe4m9bLdhFUA9LQTMMNd
Hx2v6oqXeZJTWO3yST/A+YZ+n+5GpnECt/iyZmF5+90nmP/CfRRqurmv32BbFM9P/osWwMgYGoNa
7PVLwqt8csMbRd/8TG9ZJDuwHfJtbbDaD+jG3p2CH5TcmhVRBKOHfOyKlInnQI/k9WLKUkPan5g4
0bR+vn1cyB3vQoJTpoZGw9xFxu/K0hIlJ1VbnrXtX9SVrGLcdvN7RJS8eCaFsMxHK9COidclONb1
rwG2EifmYvtXyrBFlR2U13ruPl7gzgZEADxxJwc4JtC5B9oo4Gobx029Nihv9MC2nI8G5JhSrp7Z
xkx1z86gOxNdr1OBfV8Wie2A0XfGjWPkyhCFGmcsnhtJRWnl5ui3bX+hUYe9sKTsYPPqc6EBeRiL
alyFDp3Ill12PdayA3U2h+V4iMKiSYhm4wyPTazuzuzgzHyCwSVIruCv6M05/5IgPNgvVzPn2ASY
YmL7y9EOS6dO/4VDnp0rS4F6ENiFAU3QAU4+3hh2io/76hAi3cUxPFMqof6nBIwlDTt+Pjlk6Cx+
0vS0eQgQS67qDuL7d5X4khpaq6gqVKi3YgygRSQpHxqh6NgXDwnDhqL924ks3oMzXTKsUrp/4Io5
zW6HzQ2HiDzai/4x7yYDjzj90yszT7uD5NdAti77lwDLUu2yXboS+REXz4U+VreQw/+UO924EEpX
/XaKU8QoRjA2vV0G7GS/jq38HYHanlJRf2l1j6r0Dxt2q8/mwMOwgKC2o6rSlEglO9efBMK6lIwO
2XCsfAbB9uauD9pXTQTPP5cZ+sch+BolH0YyrM4600/hKZ9ttAlOrNbkLZ/jMk41YPm6Wnx8ICOc
6vmIxSapfV3WgFBXaIZGRZ5jgYIjtSo7vI9pFB3zgD65ZzTL7n+ivgBGMC6XNUSA+LzyJ2pHJuvz
zbJdYMyWM53x//p0ttZHeE8jLb57q6F3hKLE2Ut1L4iC/EbrKpslIxZYEiw/KJWUlxjvoP/n1BX9
AfXPBwKizNOh9kfZCtgENfPZznzqwyzYB2JlHh3WLf43gPPAtSavyEY8et42WNOb+06C+54oHtle
XHdVlAQwBUGh3cGwDmbuzJDW5G0U1r0ux3Jp3SJ3l/l+gMmjXkoZZ6L30UdMty/MpxJP1COVYKIZ
l7u/VPoxOXVDhlvnnaVhn3L0YIebQSduI626XwLnDOOxv+mJXj9zdUjl3kLx02C5NU/aqg1P6lH0
tMZNjtkqGzjlgPjOUE3UMUgaaZPU9PH4JvNGsGpMeagUViJf+GBIbg5VKSi97vl5DloiUYGGiycj
63toCDmWp0M1xQD+HY/Vq+htAqpBxmWHs/lvCt0ECxIR2/i15tU5q+/kuxs119r4im0QNCZ667Mf
+pesGDGc5zq9YVemsdFwQxhVNojPbVU/u9WoNrErqGgg+cWmbmH5rmXEmh8w4YlQ1NM51moD8HkW
RNQKVyFz6hnjJzD7MLvHW7fi8D+RemxBOaFcrWpT9phHXiK1PYFuPWBZld34FP7ytIwpN4n7gB9+
ZvqyY0M9zdh14+fUMjXvFFXBRgxub7/Eo2NkUjG/9XUj//BaeQc8F12EtEWhYxfGygJ55+linaa1
jYFhC6JXJ8M2B0FxT4pf3KaeApOVmanjl8sKVQoLTx1l/oEmR/Mf1IURc20/H+PwTStdJvP6cAkg
bHcwL5NZGN+HwOEjmBJUdWet3s9kz98NTYXi585R8UEtLFvIXJQ1kAh1D6MeFpO+DmJEK8BJH9Eu
wnIi9JDBFkp1yzYf16K5SnLnaX16T3JeAs0AbXrLGeyBOKPs5zJNqqh0zwnPo3AoXxrchYFfEXEr
UOQXflpYWM+jCxYOg0ALWQYckTUmzdjRgeW2+p9R9ViBgbz7Rc2ZL3Be65OlwSZpy8JFTLjvLj5k
qyiLhdDOoIDHfmuw7YHAElA1/Kh6KhLOfYOgDRkflLrc/C7QWk3QOt8umGke+4zuHFP8lKktK6lj
Yf3OaHEJnAI0FkE1S80t5SXJIS4eAlmFhh1LxlpQVo9D+jmA9b0sm9Px8FtS5RbPcLcZwsfXuH7w
+BCSWi1Cb/VZRyAwBYpD/3pxThDE6zbqfPz1KJgHz58bNBmDKuimhp+yVDfTsqrEBYCJYkI5kQYG
J0iA0YHeguAlYWB/4dXSBW1TcvjA2q8pFz/ND5sn0+vDC8p7E73L4fctDMuw+X344UDsTDOKGlRB
qZ0Qs3MFcvcQVHOhjfzARAjo6WXLSG09yvSC50jN+GAIhfRPKGFRUCOvpoS35K8NmhNgwZYip2eu
J4YsvC5+P4tvmLsPr8JQEQ25OndUE+fZoKJ0kp4ll8f7Liq3FOjWP7VPv68cFLqYqnp8taO0nQjB
EL4L+o/Yy+yf0ksc+MMs49Jbdvq3G7zwY8PA3Iq9G7RA12jzN4wvCxfdkp6CrjI/6OROfyVCa52F
r7pmRi1+0RC598uJXs+aP9+JcpAgO23DpHF2pEPja+6BuZ91mgffudgh7w++jdhqDoChrt7+fi3m
/SQwbMq4R/sEfM+SyjIh3W8IHzQUCuFgW+6yFMflclXgbe/W7fCZmn0raje9GddAFo5AgwTPgCrv
R1KQ9KGPlI5rSOUYS8Sj5Gn3Lx58cTmj6Y1ljsFgkVjZfwCdpn1ZPiKtwSCe2PC+UAcMqWVGV8iM
Aagmy64bo4UJ3mEY9JfTeoTPFrdrRP0/IWlw43WLwlye/jAozi9IkIwXfmuc7X47dGqTcKeE/5eT
TAq3KasPoiugWRIp+1Jf2VLAYiZgagVsTC5bZJ/Y/YOii4MrzN5JzhaPQEfrudSEQT/llzUBTpRI
XoGM9KcgsgYHfOQh2c9AYSFfzWtA0gkMveCJlq9goblAPhSth5Kn+OlAlRsTV73i6JVTjKQNO3Ag
Wk69I0bVCR67La4LCzcbcgrPPER3ZOWTBVRYAuLWsKStoHOJW1VzKANW6gasY+jWwG2UC0HNiVd4
ZNwCQkRiCHnlCngzAUBwl6VHlzAdMGFyTCVmF4v0P6xN8MdB9uzA6XkTBZZibtwUWMtMI7rXgv05
Prj62Bz9z439ThBkwxkb2UrgV/akhfDZSMYAvyiERdiaKWUx39LSbxLU3PMOqCLuM538t9Br9BPd
hM8r6CENyQnya7U60/ZtnZ0FTKGS3Xl5UakyFwh741Upus0tpbSbDoJCnCOpEX+iq5tmxdh20xmZ
zOqrYvdJYT8IrIaFOUcGejJG2+PGk7Z7wqya4o2Ov/tCUbCmzuNw8J1YFd+08m45ZsDWtQYIa2Fw
1+X/77dPnrzaY/K6di5jjHI1pfucyJIx8SSjBMoITx7I/NzftQ+9lCWebNszUVFjRwgfrqgFSZP3
Zc1xAp1pmuXjDZkkmDtBM+M9AP9S7OCc81tlOV2bXc/IAnkCZsXrDBc8/82zYRVatK+uxkEkEMr5
ELGBlAKF1JbGtYFZLh/40MPpu2K1T03+MPUbUr9Vftlhd6RufGBVsBnPD/4O/n4JPh0EThhxp1LK
AKSSJrdVTwsT8dyG8IHZaQOoQLMgzdwO4HwDibnOsx2G3br2I4qV4FFS+yvMKcnijJfFzG+Ycjyc
v3lDMdVy3a02o2pKvNflx5nVeayU+AlmWLFwWjrIUnbKoteA5sE+Fdc9jQfsFTacxaAGy9ishr0r
BdjsO3rwwrECidEnGGvJMYbQbYX2FCTtMelHU9HbB6Spcw0yh5fN9+WUXJmNt3EsTBgOneiEQzLO
3YiVLcBEnP0on3gCcOB9a44vjxrKomjnhbK6JD7XM1IZERwGnGmf8Vqr4AUlZwTFstlICU2XL3Ax
fG7TVNf5ZnsDlko7V5cTTczCd3pGfpkMcOdCZGt2xAuFuOTjZuwMN4y1DtSEON18kLPf6TzK7nZ2
A9BD6DeZmO0wv8nQ9ONGSfkE6Qc4rTBEgAt4vA5GZmkbGZelh9w/CtHrWbn+ybEhpgEs1wC4et+g
Muv/AiirI+41Lf4yfGbIdwj/hYdqYnvWnK6SGkHJP5KGXo+NmKC1ptK4GVPkXkdu4boj/geZmJdj
c21KLzOfB6zAzv8tqI9WAZKaMB/9oHW9MkH2Dqi12FMusLYN6MbHHrcAuCwwynfUTYxfQeVgk6mx
nZqgcSA3sLIqHdFdtulkBLmD0zkRiLLWFgQVQrRE6cUejlqzjafGetQlYcuXmIzcMGgVb2yDXBDm
7c9MXm0zBhetcuAtN4HSgvAZ4DHKFD38wsNvYa50qzdDqBbJP9/Q5xBJKw2DOvnus1CEriXw+kd9
SzQJE5uYCib3sZqMf3AvExn1Ji9Q+btHYCM+dO+8fR09BZQ6T75irbcfXjbdw+xl+8Ne91Wiw11k
UtKoOfz5mCTJ9EYaxYqB8DapICeiJjeJ97VFsu1E1KLNy8943Bdy2CORDVFvo/w39SQu78ktqJaa
+9vyqxj8r3GlOL3KO9HcMjOYfqy+eeiOplpCpLpTSU7yXw6ErjM52sontq1ZLluhTbtnVufoYFMc
DbHFsamQBWUIE/3H7HPdZYJ9YnaIu3qMqFxcuHjAEtU7ruOeJPFEuilWo0jjc9pjGLrDZfMnGx4m
rn7JtQH11gLoBN2BVXde9Za1W6JRxYkUR6E55wchIFsomvWEqwK0lDFt80rEHvSp4AfQflHciJKZ
zm0rbqeA+fGaNAGowYaOknPcTo2/BviTPMfK4QpHf9ThDz5EUSFZFBYDpNXzCEqSwUzUQpU2z5Ft
goJhisdD4bUShBVh1WbtP8pML9Un14GBL6D8P7ZHhQ4q0ikDLnvzaMd14LhizGoe6G0khZKc2Mhk
MXU5BsEZGmtEty/YhOEt3pHMbKPyvGzv28bZpsfXG/srUKJloFfUJqWW5OZjebjV7UEW6c2eyC5z
VfvU4Ce2Apk+SMkJMBXUKOD+HSn7AHwOJiuxplhZAPXWAwlFa5KaFFFguB5XZwIkLVi1jNS2RaJJ
pbgWzRDqnxTKV55Cv11a+1a7FK8wLa447HOPPRdatjORIRGo/hmMQ+5eEI21PgRMBt4CbN2epbYs
5krAJmyfTjkuGuq++DuniebuEoJymog9kH1lxTqEcRTQoAXvHCL2BWs0wjQuZBnE54tRQLcZwDct
GDk/EGH1lkjGioALkDdH0F7vYJjGfXdfzpNudOumM8Qv4MXonXY2+5T/uln+0cYLfgxA94g+xrZK
R78bQeVkg4NUK4KCEyDstUyt3X1+bB1BA9lf9Jjmwu+EL1X2e5wTJiSJBmTxUkdDEKLWLL8cHzsx
mvU8AjviW8So8VaEGz9zphviuMve0Xrd1bACFQIfmqZDxpvn5pN7wsxWkVYd51djedrfBHGiDZWG
1/D0+rPZcKUqbTKe4X9VtKR9ds7sN5a5AvpZIjzc8lW2flaBhGRRgSlUx/1d1L2JMUCxTn2YLhvz
wQOeDWwK+P4CLvzcGViqtX+WLBLGCVt4iQ8ffEL0Hfsd8AV3MLAZgXqqK4KFjXJLEVL/c3OGedSf
NJ7ZzjMrwHMc2PsMb/R0voE8czsO3sXIAn9wC15z4ymQm7N6V5XU3R1exaM50Gt2WnGs6mlHW/yB
51v+Ec1OSSlwF9S+T679aseYk2echKZonbQN13H2UFcV4GzmKZVV3bqB/buzq+kxaxhTuMxy+5wn
4m8utNuQ6cBSbBBKN+jy+zPZumx8zA9P4r1uCCIDZ5k/S1TMPL0ZwBpMUcPUkgwxNRPskU4wSYjw
eWicD+4/C/VpY+etSYQbQDveRtz0LCPAGAtYpLXtHFTKR+kOeU2whsRmM9c0vIQ7xJXSktjqhpEp
RK3OjShTLgFM4yAsbqMQz7z1SuYremq282HA1ykbB4VAx00zUyB1PZuVZifyOgH7plfgNoMkggMP
tPY6W4fyl7KnyUGJPNuMkJqY3OP/f1AFkfXNvf8EvF2AzqQ5Vx/8F5IPNQbLKKMHeD/717CVRV1V
WUsUjzb4oJz3U9iOBTFiDh8QDqyVNuE8YPp2chfVITz6bfXRRC+16GjBfTFNUx76IEBDsWWxu477
xqw7fUyhJVTUXl6FL5oGf8M2ap5pAfRdcYoEQHwQ2+VIYBlegJPYTZsczqHWu1eDtFiKHdM1QPDk
BZht5hBwq3rumMTKlMKnI3U8VsBAug+b8+3HnpI5MAo3yxEhrDNSHRhMkNTJyfOrZFyTOGSL4EGO
MdYHhEgD5HNrPKuB4+ELUAqw9KboapvCLUIsKDQK7LFZO1EeJpBMhvfF04LDAzfsltPNdIskSLys
8Hji3wL/jZylzkQTs5n7NpDo5kF3E9CRsS37i3+PWEHU9pHCl8XY7oz+BVQAs7rN4DFN43gjJXj8
LNAmCRsryHWNEXdbK1op7ogwNYq+DCgeawtUFcslWfYuRxucTYso98Pa7fvdtFD8N2/D3JqfXQsD
BlJf5IEtf8uAm+RRZ6SSgQnbSWOo6qxppYn2cEFLgqNqHfD1n8uo2STYfL9KuScmksYkZEEvOVCO
B/qpjwlxXFh0gO+9leRzsOhznw4nDleH/0vkvdS7cb85QmxMYWB5bLQgi3L18h/PFsazQphENWXc
RodO5p/B7GJggVLWF5dHGUu5H0Q24cdvj2iZPosorWmOF6qQKX+HiYsO16/YCaKjq3Sg0l0ZamO6
4eXdSuyQv4aYCp4tzqzhaZKpbmMzoGCCxrgAFa/sRVUuWq+2FKC6m1ocnKC2wnqWdS059Q7/BPgM
u/VNLY7XuFcgorROF7hTUr/OYPYD2393zZI2+40U445fWuboX2uQtFsntXKv9dKzCE6zR20ivN75
Z44/e0KLQNu6AsISa1U61or3ELmXX7Akc55OHYoAze852jM4ijNvL9XhgLRMCiqQe1f9363wz1G1
x6jEZdsAPk6nfHR5lTNjJZ8GJc+Lkp64hyNVkfK4rk39nCoFCOrgEVZwZpfcY/Z6JQVlWKI2dPt3
ib/Y91o6ioqmA0Cs+oyjKMCw77jf01Sso87rKWF96enWHDNdJ3y3yNHN8K7+nl3+b9H4NFprKh/3
co5rNTs4PpBzQWp/hunEO+E2U7pP4Obl86yVs8m11rSyjTx0O24NXyrLK1bGGjxB9NmvQXFVoDRX
hvBtvH7sYQXwBW1XaNKz+20xCL6lIaRlP7UFWdFXIZx5UablT1PCfVv9n4b9gGjhZ4bgGxZcqv2o
GACI7M43K2+EP+zA/K7Z9S2OEXOCdsvMMS88ivT5nENWSXzY6ZVQtmGDPUsoa5BoarIn+HaxQ8pV
r8G9S+4UsxzG8jy/uQ1tx03lWxNu+s2E+C1OxbMlTB1azZkVehVazQ7l+szJc9XusHKdx0gH3CTd
/ZOGLCCgn770PplE50oUimwTw2pmVJnLxfiBGWL7m0H/tGqkHUmcnIKMvcq7R0AMdpg4pRrSMd6G
7J1oM9yiz3P5JkOXkSwUGRynRFjv8CeYNQfSHJZzIh3bSdYBIIlt0Xrz983uHNt1Hb0b/pcTjruG
N7w5Z72s2VfSNKn1XFrtMWC/mCtT6YN7NdCKbmy8+ROtSINXShLwKuLypeU+wOwOgHkYb8+aI2rO
GPcp77SBa6xq7e+MjFJaah0OaLD2hyuirK+MJmePcgl/HRKxKQfdrMRMXUanzD6tylgznzT+3H6C
iUB4DUeMiq41RMfSYpx2CoAuIj4V+6mytgNBFFIqV/K4tBzs1TCXLqExJ2kc1Fk2mu8leUMjQb//
ydhC1ZKMJq2kgnnlkxhSGT+ZP/AB4W3Edo0KTRZuAmUQpYypeKLBrFPelBVsxYhCB9Qeilly6/JW
nFbVwWt90ngIH0vA4XpuhwVzjC6nfPlB67ydaqWb4t+wsHEvxZzCell2AkT0k3cGRwXE+Q+b0f4E
d9NS8pUQwCm7fNLOtaDT+FFtLd6+XwSMXBT41F76Hu4In99Ce4CNXn0ypJnwO1TgJJooUmIih3zd
QHPZyltjX2FmU8lkCdKVWtuE40r0PL+0l7yf58jWtNF5dhxRg9k+Zx5YLLu3+PSUu8PSKt1hisAJ
bYQxrEAGztf/iIsofQmzcENS7jS2GLk0GMQQTRjbn8XTRCuQB5iUwbtoXwd5M4zSigtpzssnzQ80
UhGf8I0IEz+JnK+k6inuD6GlTI2f3SuH4zb67+TbELDOIxh7JhVuoggybiyaAqOgS5EO4/0JUucV
M2u8FHjXhTM2CW/XuUtumQm9mLDPZtOTqCUUeD3iZXS08N+y3mikRKZhHP/aPQ49rvWSf3w6NNYz
umy7uihl+31+wQksJdew6omxwcHVtl9wGUWD4sDmySn2Z+m1uY8yi4AscnhnHtQxZXrP7sr856AP
d/JUbUh9OQd9OBp4K2NvZnLzpyn/HmHBFXktxZqP5uOli/aPiPKtSpB0ZXy2V570moitYlAMsHmq
GHkAFKSpm3KKxy8eMpcGcbpQeHquIiTBdTgvfHbxORncB75WScuRg+6/yFVl/uRTxjsd9FkNlyjB
JwEr4BpeoQCT9xJX+T6TNkVbyH7wEqFJh1ZJKK8M+X727xKgYIuQz4VZ9210w+h1ufBeqLEvxKG/
xdLw0lAig+LUBJhaf67RueDpvpiDbWpQ7ah8igmSDkfPPyYI7iFamqzjskADkHuGy1azYbHs8sd6
UKAfypsqe6Mk9BkdGmClWpRo+B7GYVWVos0dgsrOVdtsjtTHJQgb02u22yXdNrntF2Bf/9OtxX6Y
ICfgBht/LEqlphyWJu5OBPrFAwZ6QJPmNa6nzWZW5jjv8QjNNV/kWTvW5H5rj04McQoBuSEassi1
9JLLI8LMgVOWTxo+ITQQZAjAPQR23YB3JthkcK4glmCRaoz86+UEZOsIPfyB4kBG9J5yTN32WeYu
+kylZFEH2zGms3Cyc76xwtXWR0WxnaqU6HLa24J6VTazXTLCYRki5OZysPR4fNZWaD0u5JE3j3/X
w+sLeJ3TG2NChL+mIWNp7XOByohYGHP2Aek6wH2MLDh0QhJdQPrRykt2xRhx8uP/DGnvkhTe/vDe
4YBcW/W2heII+ejES3q3+384enbkG99czVCSqpBkSJM1dO1Rg43sg0kNOKuJqb0Ca4uHQ8NSCbbO
mINlV9IgfXO00AcfxW+7pUGYl5fQARzYB96gRhcJJCeXGMffEhr3a0llXvjjSGbeCQlPu4dqzOXR
/x7yL59CukiUpacfpRAjqmjiMRfiA5UR/qJIIjYPXck3ENV12VQ6j87P4Og4BujR5PuhUY0rahFO
s6PfLA1phyPa72adHt3MCdoscDxaMYvlxCV82QhVHe6wqVhgzDIG/5cVx4HgbY5glDxb4mMyaewp
a+jxfovpjYWNS52T/8DhnqJgMtGqbPW/RddyiTrK+HaGs3GKYCmwfc6LCPVKiLurOfHYklloi62m
sKgm9jLl67RP+boyNKtNY+Icq2GtpEtkPcC8nhMCbcrfmEa4686ZdAEgu5+WLzMTvcY+ZzC05OHd
OVJOmPx97grkrugdwnr6w9PIP4GAaip28oL5nXk+cgd0CWciNwcnT+e4Xoha54XTQtv3cxyTuF5x
WVuHpTiCvsFV0w3S+yBNs1ZJ+ryveTie8Tc19t36NVyx8Uy3IUy/6r8lUpgu+NGobHaDJFJIznNg
mtUAmUN+M2zd7WO50SpKfEaKHUdC6qukG3W4uT5uq4NDAyjQ6+iktVyookpqoGgzmuoVhixtAxJM
y+CoKqtVxXrQ2Vi8gq/BSLeBVsEkjP+pKV8u+r18FcaUVFX1uVwvQZo255zLl5IG8nA4QW3M19Ft
s3IFtKBv4XskGCZ6CSqkTHV6r9EVfOBAYVd3AaLcTR0aznV/nPPXeba/Km1xxk5033SzqLvkM4Kk
tGkYEcpIoXyqVBoJidpAiJ8VvEwfK5jh9DCsk3BqmP5c68UAsPsFrHRWXtvX8e7RGGI98lCF6qmL
daDFuxxy44j7HZiU7vD3N9uTFZ1GnMgVdGe926A96RBMIX4CJJDDAZV4Q9SW3ggxhZRNo3mz9k5W
9iE8XwTVSUdZIMTeG8JkQ8d8zCuIevj6wJhdxhvM5yHVgE7MgJqlqOaxyfcVQPvDZbdQri9yzDQW
c1GYvd0EBp6lTqbE5bFpXMVRVgoshXt6X6Pzp90DMVLOiOuB9xwGV8E98J3KXQ+B/XXliASfrW8p
xB4w9ZXV4PQHPUC4wsAnZPpWzKDuhgghBBmdQx7rDDZafRQbIFXwF6qiGzhutHJAlGqX1wgD2f2J
fmIRH/YmOXszXsks3mXycP/vSkxeVMIF1CZ6Pey5duJ/WkU+ZDDsPWI0j3FhAqigKH97AzbRrpLk
vdFcn17NfVS6moa1Zxdh7UQF7CMYE1wsMHnUQcK5WWKHSHTlaRG1tnXZleCOGNdULM+aAQT9yC0Q
SYV/PlzHgSjP3HynDjZjwW818iUot1qFzkSWASfh6LGYuMz0ovYZLsMmWdJV1CqC9LZR9lgmJ1pq
UhwDbEFsOv258vB6CssKqXipGZyZwSXNOetrxlM7TaLyMn9inkjUkBcszbVOPocyY7IOIR9kbTru
WEPcsBYty/jSGY6t44bKcQ5sohkxYi+snDWKQzEGQtneNU2vkuWtHkl3pubPhJRxGSOW5C00cK/5
wbEV+i0HmgYJmPhOWrE5kjD9lMINFj0yv+vWcSJX1oaNhyKc5v+yAP2fCT5dh0or9Av8rPOT5V0r
002Tqp7rjDuTE09avK+rxTo/K/WUl84HpxK8bp4fHfRpEMvf5ORgYFkCsNqiPpVRLc1dTEjTxrTa
N/R+aAECpRQoZkuGNbIAzU30UFO+8Ajc1lrpynepBkLDbHWMtOzU3pvIO1cRlPZ62M8NeVAYQGGC
SI0Gbr+V4MUDOpwkfcZr0+04xeEPpU0WrN/iK2mxjwkpJDSMFmO/9PmMCXdUY3PspEZ2hhvLCQNq
X630P4p65gWO2wvYoL2EA4x2gAPxwBscLRFaWMacpJMo7C7H0bYl0L2Mk5eIU47vYDtPCtLmYols
XPRz7yMBjtzhWM/UrBKjv2voS5j1th7bvpbYRucMiunAZSuCtwdY50rHzEKYfGL2orPir0TNz+Vd
IDKmE8xAMLbRgKNU41qylXdQB1F4tfYLP9+IB4IkC6g9iqLg7vttg09xB51lcjykw/FVZQkqJS2b
S4OK9JC2fJVF0zI80v5nyMmUnSqEn6wzwddM0xEKcvEqBpGOhSn9XNFuL2pxwcpyjN6S4Dtpue4d
5mpahrGy39VBRbqIwH2uvQ6VfjAUZcnBu0zDNXkfnXNfEA23GkhnTeTLI7m4qxVaGapzVIjubiOf
UWUw0h2RBJxIC7pzmwMLoRU5JgRuBFzDcusvFLgeWKtAYwkG+egetJ/71VgztCder3apqtlSvu5v
t/2wsqOvqItYTn3wJuo90Szi7j5yDWzTQoMaz9RSyE4N6z2yT7cElqyw1FGxiQuKX9d12W89SeyE
mvu5fG9p7g3Hb1nYDSfqyF3Tq/c+wQbsfFsAhVmjxYteZy7AVJPoV44CdZraRs797FqBD/WY+Vj/
bhuHcHkIZ9svNQ4cbcdS428xv3ArfeAWR68dwAhdBMKQOd0oZl7Drp8N12OuBbG62x09SWrSK7sM
ZhdhjE7kt1zmSCVntG0Kn/p2xlxy0zGMsRy5Zqw3yqHgPnq2mjWmH2d0RAwcaoNiGSMesAXAF1Wm
kR/ofAndbNpCF0hysLqUtcjIQYh0uRNkYXOhHmHlWtxLSGv4wH9JZVEB0uTshd+pMPxV3qsNGRsJ
suntHeDmgS1Gpk97C5+4dFlzJzpkPBMRT0wGe7bF6p+LvnJQM0/lsS8e/RVn45u4z56LvPyJNPID
qdq5Pdr23heQp3fhhkFT+KQ3y941oMpBzjTHuPrgzTyM7BZ1GygAbS7pdmeabyZ5g0mPO8BomXXk
AZjylLnKay2n1QcnZA/dZnS158BjbaunpwLn/n0KhXQk2xvw7A5pOMvLAx+LqEj6b0Vq7jYMrZN5
oAZ+RNU0q362KomgFDMpIFyBfZDGr/vxPTGKAz573XSvztvj7AAdLTqYyHT27VlYEpQklDVzTKHs
5iuisUfs+DDLDPVmvpabtXa3d42oKK+naF117lYw3CU+a7zrP1j6L7o6zPk+7MZcpX4Vqb5Oc8Fi
Sko1i4VMUmB8iZH1O/QEc5m03nV7YwSmWhb/EU5U8/cyE4NHYRxzJCMml9PFKEnmZN+/9NnSrxJp
QIiiG5vNiCI1uSokAFRiv6o8heJFmMYX8s/XW5n8yvOsaBdAiN22JCV6Y6eU2kF7ENJj8ycVrXtc
GhYSJrnESZiQlePbx1h4IcHGASWI7/QI2ENl9b4vxKGVs6eezOD5NFrpxuHdXeiV2INCgaP4HYo5
kpaawg5JiQgPsI1FfK4qXYlSWMgoJ2Zg2dcERXzjrGqrUW5rliW72P6+/uH3wMtO39WoMl5MrfLD
cdDE4LlKNz6092lYHU9vwzgM+2c3Y2WtN6n3npInutYZz2rUGOkt+0gMbr0UROdaQNG0no/KFzp5
zVUsr6eyI2P6V+tZD7W6633emtTMJrVQF+7MMxjEbX3I359A/Zg3rXwYcqTlf7COcYmM7vSfyyDZ
2mb56r4vSgD0LFy7pixEGv/yaoeMmYuFJzrdagBFs24IhmY7SPFEzt6+qm57OaroWEY8dnohHgFy
D1b7zKT984dtD+SJ8aQ3/Xg8OtDLy/PXK70Td4jHJ4XaZFWLWWqUSxxkjd7L4+6ggaOrsy1Cf+VB
QeC79RhYA16dWvereJHFP9kG00cufY8C4Z/Mh0BnK4M/ZEWVoEhmMJimzvMKNxoOgpwrdGT8/2+5
04PmhoWANeSk0OkQgQxYX3K6A4eB2dTkpcOROomvJX4WqMFKAjbS3Vn0xnv8dp/epxEss83T5HVj
pscBYCDqUQy0l1vdaEOBHlv1DaiMob+rgMRAoUgi0zE3WLQziQYAvlZglARDFlSxpfre1PlB0k/7
E1wCglkM5i3E2Gs4D4c1PWSV9KizfdmtKxbeu8ue9EeK/WRol+wqAKDuIBID+vMYdcPNwsq0tglT
EKtDF4hQxWbrF9FuW3GiWzZGS/65HwvZLuV12+6bDYDuaS1qot4W4opfmND09VlvjsZpVhCwASsx
Ee/7HJfJpwj41rrW5apHhdW69z0b7Ef6ls8KWhGNRXS1j+9oNs9qpBK0Z2T5632SOvpxG71ikSpI
gcjp65yiLsMT8sCucmmYvR5mbesKwu76creGkvCm/fcuU10QUzWsSWkVXAETIZjPL5W5jCuI5NnX
CljyQY8i5vjgfstzwgzWdTXx5nIa7ccUoHUlDfO+iHURw2wIXhe+SE2cx8VZAqgH9JZ/rtg9SY2M
mIn5uB+2GtINJj7RstjC+y45LN/Km2lFCpRnxNPUYPi8rRubEaqIA/NWrkeNqDPdFfTucrw9wxgZ
DEajbMCrc9M8Dp2pSJaOMRmdk2IDJdER4TpXlH6lu8QA3h79mpmo6I6wwv8gxBPG/9+cQcyJwuZQ
HUT1OySCstep3Zhyro4RYSqLzfgbR8my2EorH/4ELQBPdWUe7C5pbvRVZnZmkypajOYS0zSHAsOx
1VIjjh+Ww1yHhyw9ABHhwKktjbZwpWWnYu9Si4umJ3FYIq+0tofDl1glUo+kP6yJYAzrxFMv5uEp
/ws5+Cn/xXmB9HM+tMo+G0Z4mlxLzYwOzcqwUb+lK4ULoTXuU1TzJquAPq/l1FOSi6cIc/FxY5AR
mx8Xr2MSxgXwsW7wfZuU4SBq/1D8IgTgB/eMa79+7VV9A2fp1DuMAc1N+h9myjCKmLLYHtM7Wr4S
m8i7NGazhKLEDxCVdwW5+B4cMo2wllNpOQnU4J92mdBfULCvbKVb3wlUTu59YxGfHKScnH0t/eh6
dRtZ3PnI8VgHjpHAnfKraNMS6GOtfkl7YE9SKJ4RdnwA1mIiAZLlYq2EI4sv8jYfSpxAc8AqQU5G
yQv4dwjUlURT+eCnD6futyQajOHuPnPUFXWL+NPyXuh6BhMRYKcRGesh7JsdYwctrx+TOBq3wwGr
Ycs46t6E7Y/4+iKZxsJIFkujje8F8k7AvQd5nAsWaq5g+A6ZNrh298jrIKQ2XiPWdx2f61a5qElL
uOkr7HA8ZNskPSwmrF4CjUC4rW3l083NW6oJt7X2jqt5VkpqAoUq0KkKL6Nri6n5ixTTuGN4xOYd
ONAY/Oq5xthMEJLWgs/MFMV20LJlqiJoG0NBm/RI5vl6oFDBeciEc9O/caN1ZUtl9BJuv/V9spnA
IuQpVu4q1pPqOt98XgVc1/QESIztozxDEQZv2k+mJTyPyws68DINdmsTdPXaAxvDwYAJQ9PtotIh
BF7r7QqSmCiCFLNg7y3b7wKYQKThWbq0R8e0SvUPPcdRLJsH/GaQKAm9VLfYe8Stte+f9uk3OFVJ
sCBw/NF6Igh91LF7cSq4R1zwf4lEXUoTy96BMpkR0orJYSvh9VAJvHVeijawSMjeaYHbjdJ0dUAy
uNOzmKawufklOj72qPvYC/jXK5iSXnQ4qYzUv1FGfkPloiR4Ay/bRcpkd3qVziRvHNztgYJsYVaz
JPwHg2adZ3rtOzyizidMZ3so0nVTdLbtwsOm1sYyMAshxTVBg6aVeAHdP6cRjs2jxPvhzKrlqKMj
+pFEaF09DJfrwraDtB1cPGNvCvoIsioVDlRm8ONeu8OaFzY+Bw32PIKWrXfnGbPJaB6ZQK4C+Fy2
F6x5uCLTDOcCBmyMCzKBHaBtQr6YPO6xYAVArZBmiQbrXXY08dK4up4+iQpohjdG8veYm9wnGlNK
F+mptwg5U+8u5Vjou7ZIBj3JrZc9vfQrJAXI/Kbr+2gTTS1KTKEU3uvoUYKtDX1cIBvNeMqw0ZRF
lN+7TS60zvCNuMNQUR0KKS7p2D5S0dtJ1WLZkTFpallDC1YSSrL2546WDOx64yrquS4JMJWGN7Ka
3SB72LbV4mfxHGYI3T1b926C/0JYO3qDc2qNbg0Q+dVroDRSoYFfnmYMzFAqg2s0Z0LNvhDx0s1w
XThh1q48ewjOYV1WLnqg//Ytxtp3eQbj6bS3bq/8PQIlwo+p/3a6aG9AVgKIg2frnLpZFnpo1V30
FeuZwJ0Pc5uxUXI7xKV290Yl2ykZw1w5d+F8vH1m5YzF653tOy2f0McM/67sO7cTUMpHbJrJQSaU
2qam3k7apfbuANwYXpTjJTHnHWWDlN1t7NoVORcqBonaC42d05Eb2XPWFFnASG7hLCJJO09juiEf
kQUGoqz46fDxKCvvtBUal+T++6v4nqwPP30BgFaCCCxbqaalKS/AX5gMcT3fMyUUPLdRZA+4RMnA
Jk0Wcb6GRgkYx1ta7s9kkqOb/JSAS9AngVl7Cyof3GZmk3CmZi58MhAsYoXCWGxbTeWeytZIy4nS
UkbuwMfT0lHNQZlSR+lAqBPnFEUx5rU/BHUuMn2Bl8lOeDmbDQ0np4hRUnh1zVvTptoRUN6QdrsT
YodU434+gSGjftF9PoU4RbfLCqpOpqc16zYSg6/YAze/N1Jj2lY0orF5jUkOWd+XjVGKGaxlQ/E2
oghUzdDv23HMY6UmvUaXKVaKwRMeQpxO3g4PKr4GSan6zTN76R77OOmBXCImZBlR/mpj83w6BnUA
GtNNoBwD3arrJ+3R6cjpPe8OaeZ6pbwfTE7pQUnU9cgNG+uItq+n8bKV2rM9Sw4DOL/wVKLFFar4
jbdkcJY5bdtjXw0/MJTwpGVJsOPtNWXYS87BJPDLz1IeTr3O5acngdg0wEjumfpCFUj2j51cMjcu
i1ty6XsvftCaHcKGcOiNLIJnS+/QEYERfLksx01449x1fJcCEB3cPy8xZrh5FNio0gNQ6Y58zQQ1
WGh9juJuy+tmgZ11sPuOA5jMnYT7AdzP+v18jZ0Ws48q2jVPcQW214Kia2wld43k5OtSiLcEoM3D
zka0GufIN7PNh0O6o2b3cnbWzylwnciibDIXWoWDT5cqlLUIWfrja/95timZqdIdbNSrPF89h/44
1SE4zQ7yyFH7S8Ser+z9o1qo9eVlhgmVyvtc3KvQ3C/ozxcCDMxv7NOinmaCBg17F5FMGhs42r7w
6/XvtHWJXdF1HO0A4cCSgePk2SU4/lzFwHCT13oVUKfULQpfvVcNTOY9KJyWtCuBsjvKsL2jiuIW
c8Kq1TcOwNaAPmKW8dXl2coNejm1p34pHRRJmN5XneEydAizYYvZn6O528Ka5qkivqGD4YsbVdck
//qrTvnfQJrTYXYXIY9MqztaVsaNkfF92S9o4T1kFSGk/2jBJMia2jtpFHyDDiD0l6ZBDlKYiUYy
4sxsskymQhJqNPcLR+lNeO4diXFfdpwyr7oKpcinDAOOM/4BheZCgSJ8V65/+M4ETEOIggJnKI0K
jeK8lxbU7hCIzd5uJqQqu6PdJCH2HCKaZj11LMVtUWvDkkzNlxjtetAV0IlALPEirTiAdQMZWdgP
nShrgyxnRTH6sAL5CB3RDEVSwjuEsTBlJPJ22x8Ml7D5620nddq9MyuLGnE718WmaVwNyd685khf
UqKt0KWEs1S5AA+wRC220XUZp+ISnjNZFAtKYnOwC70k2RhZINwqXGPuy5hrENH+2sXF0xRGLmoY
u+IJCDvrc6k29S/b5lw/8jk1dC+Z1IWqfYKaGOxk4c8Tv5eAb6SxoI0Ggl+WWG31BmZHTWrjXrtf
rYKVjiOZdPfaZy9DcYYcdfJVUnauBkIwyzBpv4BHPVHvF3qn4Ah6ivUVSwXi1U90/J2u/td31lyA
qsETkz0RnvMcxeJLqpcfx9shRum9wRwi8Y/YfqYRSiajVS6lxYjQu6DW+nxp+jnZk3/xwLQ3WxGX
Ovo4pWc3VYOmFeNtyEVk3/qfGREOqe/X1sIMkhmoEXfyzWm50OeLdyRCMAuVzs8tpCSnZ2mLOr82
cmZVEQGtpGp3awNmN7enUaiH5r6g5uaki02Gmi+7ZLZRoG5xh3UD7jQDbpDgUP4E877zaG0L1izI
xmJ8cQnJpYABl/ZFuecf9px23fLrrDspIExZ1G5VtB3EJNQS2mQUxCV/vGMIyWhwYFC6VqwvRs/g
QFRdW4qMVMzl+u8h8ElgEJc/RJXMatBvCE3TfsBUUTQ58ZUexxEvyHqXLf1zS9CzslHQtdq/dwTz
5fv7TMt2XxLjkt632ImGKT2E3EpXW7tZ81/c5qXzMpn4OPYyxz7zSjqV5paUjp1mE4gRZ3sRap8h
spsoOHFaeiNRmMWJ/ybksxFePkYrgX8fXLkeBm4U+gFzJOGmCcZ+E6v1x+yzX4uvLObfmXkkxjv/
n6kloXRugQM8d/nTkrtEGhBiTLirp5lUQI5sN3z3U0pLyP/9gROfGVDH2g0LtkOiVc0cIwjoud/7
XgB96fmP8Bpz6uHRZPzpSZ1FuNtsH88p2j1S8bnDLLt9p5JTeBKazp32YUwTGJDCrt94OnB3degC
DxSc5PVJ0/l2tct2hx4bNnOS14S0Eoo/zPiMP8aSwu+PbdLRdPv4goyVtkQFADXJQF2tNbid1Afh
1S/SvMzf5NsRVLvMsg1pWxn2GVqmqBNzovYsrwFVD78Z48gu795LzuWRmrs+uxPi6FMgbWCKvOqi
HM0vIe/wZrfqCztrI2InafVDPHr/XemzQ3Hka9gqrvbrjoEDFswild9uq7wDXZumLlVouaxeN/cw
OiiADadUh4Vp7jOiCyjFYYI8KgDLm3czEQ5vUjFEjrVHXxdMTDw+c03lvrbzso9H6WrQNc5TNhnW
EAJrMhOBZ0XMMnCAkSrfumT9TVsdxyO+rCmpsNhXx6F2pGqUdfSHpcFJ5sMkR6a++NI8NVH3jgxk
BNh8T5cWScgh/cUCMV4TMYdX+NvmGw3ESMO9T6nzVihjpO1/knH7TyKUg71vV32DNwXBUcdGsZPs
dfotiXPV+/xghWkF8SNgqpdzF7zUudKMgWiJTVrkLycWOjq51Pt/lOZuxcoT980qSFQJHUuBZG9C
BuMy+gkao7lcyHaTGN4mltL6cnPakTJiUWgsDGkgTF8F5tMAhzFtTZvyYDwD2HxVh8vLHrPLFXeB
vxyIJHcYwVMhpr1DMITRQgMc1krN0ue/2PIToDqG5851KkBugkWU0+yo5QwgObhQYhBRx6QgHVU7
7uPOv9LSD2FWBnxWfVtzN1+DRxI6ZaBUki2iTqOxXqxLkDCJSw5o/4dg6l2wc/HTiPwe1qWM3XXZ
zG4BZgwyq/Xb1UkkrUEd41XIbOKeHN+hgnuQ05Li/h6L80XUD9ZjuNrv7JcmXcTCOV8a3dIzoGjZ
iJxtOZVBDO14LX4U+jZ30BnS2dpTS8B6H51VnpJRIrs967zhHYCHkMSGR6Q04k/vvyW9yOzhkcyD
rPBJOpPizwKnUCDJnOfeDDr5kq5wn1oMI8UAR6r3a6fTc1PSM3dRQqKg1ThViWc951LhdH1qhYhG
alLlYCNXa9ZyYTrxYs++PZvw55Swa/CYSIFKVFHdRU2eBbodwjkJum74Z2veHK5zc6RWJlzT4cte
6yNxqVR6liUZ9S4c7KIU8AIq3iQGAYLOC4oSswOHL+7CJCvoK9i4Kh65Jh4repfM7+9gAKMfzerM
TzZG/1TtCq5+tNxhnx9LDcA0LpRPeK6SVmC/L7Ejc3w3HdeI4IirBv/7cb1/kciOqgvZxut0IcKE
QaZlnVMOrLw2V5kNq7UNdaiSZzv43dLLI+UMM+SY1KPq6E/jhpPc9mq/18hf8PMg0s0ky+xOEvsO
azKYl2RIWWYvgYJNSQnUjUT3uCqiQpHcHD4UBxwCU+4Ubg0KKzmEO4SpGEq5W9S3wVpZzxZmBzbR
2qMTEbznl07ntdP9dVXZKtVLsj7QfdRtapSUxJxmr7Opgw4tu3oFL/Xt6AJ4lv0Do1qxYc2I5nAW
iIWb/MQBEPaeuBuT5pptM420k8HVvtJITfyLKKVYOGF3MkQTnyLxoZzi6Zzt8XwzLzUjWw4ybPqM
6BXKclrNdSd8qsA4giggQRm+QIpnzUna2ql2/ZLGoeE+uC0DeA+uP93UP985EHst6o5d+bgnx2n4
n+sWLGhKn+TxwNZKMGyEhd43q981jtg5/95nRn9aeAJOEMszWkQPZIq9U0flNpIZh2fBNzCOdE2u
3XX8lhGDl8jkbvlrTYqr9GF1GvSoxWPggUQQA4jeK6BuVEruW25aC72slH3mbnen22Bn2+mOI4F5
SQ9tsbeWwmXbACyPKippMdcUPyRmmwCkrG33SDM7qC43qDOrpUY6vXcYm/xcjyjKSEPSXhn8uYLQ
ZXmQoD3dL/hu5ZYBVi8CBLWF7Z3M2yOVwDiyy5cJx4jDUsGzIZd8N526HYwQ2JEkk05xVE5DF1gT
AcbnGlcoylt++VeDrwXbxyHDBHUwp3wkuCxH4Q/02TQ8Rahn8xdSxUwr07PH+YgXJE9R/r0QHXmI
0BbtMw4lxID0ptMUflgw0EkCRqG3I+P4N+iLB3A10tvQ2WBhbmcBl14QO/hJmx4nc+w/A0EZaK1e
b6ER5FiMEqtQf3vTtd/SPCwRmIxOQmOaXY5gihb3aSyW85F1os8XgewiGhBOA5qfIrqs09qsKXc6
BPjJ/hysbB72LxLmt8ReY+OGJipE1eAnsTr/9ZMSZ77uXleCjJC2Xi/GYrGdrE1vqTL86AtQXMUc
+0Zg5B9iqs5ZFpxjJhwpjnN3MZeShu7n8PAntNNQnzvIOaLtxI4XiaawdYunHBdwV7q0ofgiyfcA
b0T0OKB3K3NAoqQ9sMLRMzZbTUlls7q+sA/hXvZ4aUv1lA+UcSzSp2/xnA6gHJIasTL59myMMVF3
W11AhQ4o0Hs7YxO2Gq8oF4O71suAyjwveGQCWa9FBzKGqEjzsSx/jLaqxgXJxMD4PM/XpcUOuI42
UpffW3jtWJmp7B9qgOuv9fO0Vx3PKZJBx3xR0JEvu5Fw+xOgJ2j+AiaGNO+lUxdEB1pX7Og44AHo
DmLb3B5oRk9OFRAHQs+5ix+fXzQ/zu/ir5K7LH2M2+D0UeiTLd6FMiyCWFB3AZPcQQiMq2z5c58y
Vf0t/xZBIqB0w3ClPtqaZIDToRBRi/yqy+5i03xku18NhrZfQKO7uHa5AcNn49UD+tuKLoD3QvT8
9oBflPPYJie2dX3LTywizT3luP6cyFUjlYXgK7RXYhP1b7wAmC+S+VlJ5abxdr7CStZB9b9LmaEL
/Sa8dKfSFXsvDxLMOz2zawWXHC8pTqXT2FR+eE4P4+ZKNmajuoYOPkZdG+2BSp7vYSZzs8Kgp8NN
Irw8oXMQWM1asCnAN9hSmIKI1CMsSvbp+ES+b5M+8y26x2GvwjV2gAL2iPXOJ2l2SoXMZ6idOkJv
Z/bcLRyKDm3MBKxnbAlKEM886jiovMrlif6fzMvS0XGw9xr+yfUqgwBiPlLC+3vpUrcjiiUS1PLi
NIMIPUI4qH9x5jK674Q4MQRSJoV68BFruZv7Aq8sPVR7PBbEL/KR9asBk0DL/a3/LoASoOVsee/9
r1eYF9mdg3yvcqNzC0hWgDPRx+FQ5i9GYDZFxq5oJEf62h6DJhG36A86urcrfnVAm1ayHpwlZGqS
OfTtvxGdvJMA5JJECnR5RFsKTqmSZk97uqR2Pja4pbw5JSCZJpJghr31wTXQJOWUIHmxVOv95whL
kKPLBVIsJb1O8G1z7SVsfsfvQZWF3GaQqhxU8i5ih+u2k5P4aF2Y3QovOp3PGqY/Nk/PTspheAlU
gksvwjrAc1ap/xeu+ZRPaIUS3kqvlTZTSO2RT+HVY2fjNhzllTvqccbxxKzrU3unssX8mlQJsG55
am4a2A1fIl5Cao1zqVlkvxuB8vjYKntXCq/PxO37wcpP/2meklgOsOeYnxLl/aExOiRovITz/qbj
ycsc3D6/lhbgwa+OKxQX12qtzSKqV/cGyZtlpJ3T4IeuhUEIyqfLty/BfYBFl+l4rCNmX0RyVAGj
ywyKVyZ23FUXlLII8QRn7KpBG1iFANZhH0vY+rAOrYdRA0JpidMjKecsagasHFN9r+FbkkcOmyJ2
f6S4sqwQnKkzS9EawyFsCPPk8GoyRiOWi6oktrO83ySwhp157oVEFNxA9CAZwWCfCmayQFT3auc5
S8hc+34KOvlBqrSB85icNuja7Y6cLYBXBeedVMJWzotnzIE2OOMuomNHNIwq8d8x+uM3HrOJTw9Y
cgXuwnHCuwPqQdJqwfenW5c3LKSmpLGL0WLXDDyyOO0gR0eF5O5gAnP+MUPpxiWMlV0ITERDMm27
rDYVOnE1JSlWsYhF57FcXVvioH5RW17dCZk+vjy4JwXNOkXoU6Ah6E0t5BPNfa37Pqcxfuuwwn95
xeeMsAqmxijo2ksF7VMM6piqXuqOMradcT0qPRAMG2Up/mF0rwyxwDEHtYgbRbjcshzQSdd+es9q
j3Jwr/MxjfGM7cFy5xeIZMojbq5yYB0U5lBaib7DWxCLf+BOBPV65zvr2QSn1NPjXAU5U5e9w/PB
S3AyEVJr9JP2wZfGgqLTyvDJpAm9RH+14GYSMu0e+s7TSzvUg/PFPc+4MHl9rBwsewtZEvhX+IET
JfU/T24e701HguX+fN/UROvmUm90i2eAciWJAk9z074eMEpar8CK57+er0LoZB4/kXv/+1b4eyRx
ejz4rWCGisWuvHpVdXhSUGauEecPK3Q68DC2uSVS/fTMRiM7yvbQY6DwOHhTM9MdbcJ5gc+xaNN8
YSYpGh+9yVk6DOSl4XYN8VQ4raeHejCnrgKgosSaNnedmV/VWc4A1JPgne27m+E5sfj1W19AE01V
FquwpuZjVY/aC0grMgmYH4TrFodCjD8svMYM5tZJkbvudfunc9jo1yNgFiiAAn5KsAiKJZ20Nb9q
jEhy2yXIQPyQyDRM6IAgWbV44NGZ8eQ2EgJoJ8QeddPpF8D7Sw/dghRYwXmkM7E7Q2gorNaQ0v02
Ph0fX/0ZVab984BiITVEF0FQliQeOJyk38jciHFqHWqQfHhBntgdLuCpyBWIX0NprA0Zc7ciTBGP
WUjBLg9RRwnwcym0Yz4An6Th19P3GdPATbk4t+EvVFwcOtjsQ+i1eUQFVuxFm14GH2F+/QUx/qBP
st52bMJt8K5C7giqYCYWM83bhVm5MvOJdC1gbG0hpany1PiEnS/ugNllt6LMUgWcY/m4rYxvXQxB
ulaWzHL+b0a/RICUWrEfMy2nWRnZ0b4ZCqJ71c/zXyyOQTwB9hVFDp7mnXWkFHBkGDLJ5N5XLvVo
1iS8xkooisVexOizPP7wg9IUYuYFNLWgIB+y2Oaw5JraeZ7PZDcEE4NYK4plgk17QawWJNig9V+r
cna6xWIpW8R46aZCOJN/Ncj6f2Y5wxfx8FBfLDqSbIUAlfoQJhDMleGMytNRf9UAcCgfvBtSR8U6
g+KFfh8F+iFM+UdDTqgiFqbCiCB3/s0lgLztyKdhTorgyw+PCAL3XozsOHk9yxG4Nc2lS/VMYjy7
Aa3gqsnsCQ0s99I78qoKT8z5AGRAyN+z2JUHrsVhVvLNLvrEAJtfcrGk3SC9hBgkwdR93gHLLb7/
9d+uTHv6e4DgQ+BUsT9GIpAnrE4GddQZtFUV84uz+ICYTEZCH3I+BHaOUZocutR5ShHWnghedYmu
vJHx3PVUgU2qT8HFTlCidQoUtM5ZusSa9pg4f+vTLd6QpZzUO55IIAZnQcQP+drx1Bdz1cmm9+Ut
9o9dep0pbbbeinQ2NlGqwcnyYRxkzBQjU/CAaFGreZjaWN5HNYUAPjwzhE0H3JaVOYpMtP/ciJc6
vjiMVyJXhzUBYcwi61SvvunspFfne4djPwcs/tqctKKA0IVfmd/6d40FEpSdAbqFH9bBChspVK5q
Cl9K6FauJ7A0hdTkzbCNZ8L+O+KYmiALJewKoeq7mgO6OHKXdQPfw/OK1mTRy1dGo6gTcSc3eSXr
B6S6w4uso3Fi3cgw6PZ67NzVBaqcdLX0c+psYuVZsnvB/YVUpPIO8bx0NtyHV1Lw8+DvnwovjVQ4
3SsE5rrvagMQlvbrdlL+2FgYzbsfCWIF+ETDw3qUwaNU3RjA89PqfX6/UzX7uJTtMf4iw9YtbJ9E
gxYzmIolm81uCB7+InKXvocG9/IN1+63AjHfnFf530LKiGd533Bdgefikg0QundwORA2f/ZsI023
YjAq/gtcOyb3RYEV5K3W5E5vi3yeubTIda7eGxnahPPTeGpsMPSx0oIyFyhF3BGs+fGjulFLhT8w
TrSOg6Bx7L5LQuCMARzdYy/6S82q5zu+2/IIGteDtadCO16W2F5wZYkBOYBdsYyM0alik8S5WkXU
OIWDMyb5uEE0VMA9N8IoFPlXmSXgRglHgDrLn3fRhNQ4oxpnOmL3ZZGtOasqd6c8TzrT0G9i5Asy
JYByEJdKqnkzIfD0Xi2lWDV9pFCTiq5CkgJ04w+wM8oxwYqdcRX21knXv6zA0X0UMjg3wpYLXnq/
Y7jSSUiLoBStLF1aoVNNRi+Bb6csNbFAjgTJaDJS+91d2Kk4EnZlE7rlGfsw69TKZD1p7EshSh2R
K541eOqsPXtwd9snLPUlPls2lQxoAFrhSbozvy0TEHAYBm+p/XE9HQpS22wDKM303wJT4onnXHmy
40UNg6MNanaqS/XtqOvNVm+ok3OSoARG9qgOYfaWD/Gy2Xfob/FdbB5UnGrtMqCq506X25J7ztK1
9ZFRnwJ2c4yN2h71Y3Rh16ouCGyXsK6b9PaAvo3WIydElGmrqahXBDShuge9ZW+W6A4Fkz6T+Pp7
fBmKi4lDGWWJavy0gQyRQ4R4rR8hUoBpPZd/MiXXAEr89vL0NUZ5hpGPlYiN/5Av79VxIn/4DHQM
uh01XKgsxp4UI9V7V2Xe4QN7QbTHk6qgZEVPRqVWi4ZyvZe5jCFdMSk+Z7/f1J/CTUA/eEAaAP7e
rLIe7AJTcCL1CTR6E0gfISWRwPG8uD/RaNajnzgFE2kuLvI++0wZ/Zv41BN9YtNVBDYKAh8cBuyz
Y8goSNiXoYf63B/2THHQvLOpSFBvEtWJGBq7YA+wKJRGQtcKA5eSXrOryccrq+O7vbJ38oysnawl
BbYG2MdHCJhu5KbIi4q+fU1URBV7LnH8y0wVMenvwmlcZF4pYpYsxQPCHToAOaYB1tvuKQOCLhPi
QoEQn1wyjhQAfgjUxj+MKLoCfAK5waeh6NWDBkGnjMPyu2UMblUeqmUGr4Xt9flL2iEOyQh3uRKL
0nu6GiacoS3iUrh7Yvf5XoQ9kSxQ5UTrxgh4Bw/O7osLMQbPIji7NwUBagGRXzuis4fdEc/fo6Xj
Ecz9q+8Eh9ezwgzbZkGm7FXdwlEuzkDwu02jkySrrNGD8i7djuZXBaOJ4w5k0/zRpgFS7jgrty6R
rLpZBRAJ9N7ry+x9O2ia5Dsk1XVWbldcYYqAeLIpOYW1eWaQu0rXh1C1+m0z5BY3M1MoE9JP7TUo
ydjX7wIWt5US/3XwF/Z0/N5VIb1AVPXRRqDe8S8p4xbu2BO0zOQjQmv9oWy3/hBc4TCDuhoE4wMc
sdRZB3ay/3MqkhTwXw3uOxs5dSK6iXF5kv9p4VJrWV4eCgpRqGusT8xf/MS3JPPqKzVMKqang/o8
zdwfwGM74jadXWoZpL0qje1w1JoQ80OpKaDdb4/qhgoYQc2QrR/v91YbeBUK0nPjywjrHpxhKLhj
gdyr6Z6BMVeCAoWU2q/KJe3KMOGH236iQ99PsZkZ8qhYQLbEjFbGax5h7GgSIX3VPd5Abc4e+bcT
SFYYdhMq0tt8+j7p0bKYlHpFMq71L5h23XNsBxTCN8eePHq/93aHDRQKcPwijDc7JnpIfrySP2xU
Z0SAp5RhI4j+ovlkCI3gwFgXiESrTNq/Yq+ci7FGkJSia5bZjrcxHdS2yxRdhxX2WNUxtjiMqqlM
FaKZAhk40tobyG0lm0IUGQdbPRk30RtKFS9eB/hB62WnzWjw4fpHYbZJBX/WACABOW+X1UbdelgO
ATYwEAIc2awau0xGJ95ebePNp5wgpdb8/7r25CjL8I9mhcC3tmAa4084OqcWJqJHaVXfgoBswSNo
ojyg9aFO143wOaj0Rnly8IMlSqZhAXxN5U0LelzGa3R1v4okPckHdMqtucNE21FN/KZW38nbJ7df
54evVQsXXcOfe0sTxsS8jNSpxcVHXU+NXxKMuDV3Gjf3ICMi/Gtq8FD8BXUTza4KYMyb5F8Wv572
WcaMIovams3NxIKh7DZw/WHCnQdHcqj8s+FRJwvtnzBvUp7kFHR5l+TcLqC8B5hO9po9Y2DqvW1O
SzDyMph3DcyakC6Ax8Hr/619/o0WS5mtWw/1fTyn/QQ/HPhP2dP7vnWMFdJM/+nM0LUBte2Niwpp
AKuaUhOMRNrQLcj4tCfIfHwE0Xto7IXXU+2rbAulcpdKGnt7gxh87Wl+wB5JGejkX6WQVPNsYTMV
HvWnW303waKbHuUl7YPYYOQ3LuCSI0NivSqfox/gYqOopIxUaurmNI2/+0OxyWymSlslnhQFZrZo
ZUR7/dF3nxB0fa5etVOY88W28tgR9Y+SH2kx9rLlFwF8fQhZu+LgQ1Tmv2EVaMTZWgSCjK0T5CJi
j1PjIzMJuR8l3/7nnqcWH8viEkWjOvzfjparo5QykyvzaBWyKzi4eP5Xz4Ntr68lZDWbFng030f2
zyU20zfFtAt41hvjhfzha0nIuTiKZVaPBb49gdtKVRxpg1jStF/Mv8dT/eOPe6YDErlsbe8zP5A4
FBF/2RZIilW82hef9QbTve1sxn0YWFKhozjN7xg665rx3fbjnxtPzwT5NPUeJHvmqLSN5zEkgWlL
7HGO0SsuiTMRF8639/tgI8pby0Z2cQfj8mS/I/CDVVX3auoLH7M8o4sM89vh3UrMBWmsu5UyaDqE
2sxwwz/hyYVjxigO/Xny7Tqbsy/lz9TaaRSYPrRpiS+QHglOhuEAnAVXOSec+X2DbEKxM0/Y639A
WmlNYzz+MALvnSOpbylhrIAyKHwr3VgzJa6svJAurQmwG7axpBhq+8JalEFS197dSQRzcTSXDwu9
vstov73fFy7P9zCu6UbjnfNVQdMlCqmM3Bp5ZUbp87I+JYS3yHUOOV8YmVD7mFekGtxGah66KLBV
MFKCXo4aCER/QEii9UYKy/K/lO7rzrq2fkTBzSgIsobAL0763quUoiPEd8Pkh9Lwhz+5KHSjKQnf
C4Yd+UsA1ybL0oKsaV+l2s7Ib5KvgZZWBUH7UNXAsT4iRUKD1T/Srq58wTg/MekJARN1WJIuGjQs
Y6j+I7zlnBKuvtr0MMZMS8ZokP3qUtQ8OKBqP3cNRLZ1OnpYSPSE1Wr8OecjF5niknBXVN51EzNb
Ucd4MNZnpJiVvfYnN5bmLT2d2r6/Go1Z9CsXz/FK+iBGg8YGBQlBx2r7bsr2ol5ag2ATrLw3rdo3
21iqY/tjM4jZRube77zea1X3tk4pQUpz1dkZIBIYxB8NDquwBSr0RDY6jYDlI0WqTILGo34qzJIn
hPmWY9Qa3TtyK5N6EKYrCxRzx+RqMNpV9jXdEEopQo6/jHDiSyIxFcszMdQc3zP4gKIj9LGHtknt
lkomHU7AbMeC/DnKR8fBiJlqC2iTeGnCg83DCdt2irTcXykig9OHv1EVPH0NQ/GSOV0uw53AoXNH
t99QJ9iiFWVueT8bWZHIN4dHrGJ5GN7XwNop/v8TH7DFa4ijf6UtRqW8Vo2VDaFS8y/JzQDFtwa1
ISHgLwf1SRFPJGRzSWfhDiytWlRyCeJZh6yKdgV78xiXLfTvDtxN9vEBAUDiI994Q8TINQFZM/CT
FGH29VqXLgRL13NdYx2IgWAbO3TQHtkcRiCMiqCOm5s6G9wfhZR2voKuMeitBR4SGh1zmqShs9ri
/8MO82jKfVhVBP2a0dNIGPNJgK3ZE8x6R06wO00DvEjJ1mt0ZfxoURNFpMR99tqzKxsQ3f2qyk72
L33Ub7UkuMCqN2AsTZaw5VFmGgLyMBDL3lHu01gXkd15e7TLUz7a7YLq+c0rxr6LeUTUTe/QLD7V
65yocYXERCaYMK897nvipvAZQMKP73mxMt+7MUrT50UzJcLYTXhK3z/RrJEUReIicofir7pqTThk
UHT4yiKgoFBzHKdnVO4ReG99UdMuhc7k8ikXINpwtiU9m0E20c8/2hhQ5X2uBaLU3K0PVj1HPFsV
yIW56SXOmovxFeq9kA0vSG9POm6AWMn8lUbMLqloe5156LoqtE+mdGjp3wYy+xdeKARlzwdj3Xu7
jWRUHfdGxFARFm20ZFnOT3fLXIhiBxKVUEUPc4/7bYJ2K92w3T5ND4hIvkAgVWB6UTpKBHGWv/vU
Wl4ah5AIUb9LKvZ7Sp8jp48unOmZj2MVEVS+8vmlmWQ1FNby7rGIlcF8nht7QFFFmSh4c/ogDH5o
RIu+3RRMDgPMCR+1+PlRvubJ1yh2auaekMmrC4VxAyQ9EiK8aQPC5jqftgQ/VWqG7I8SOvkJEhLk
k7tZ0XwoD1F6M58NySicZijAOsEkERpsdSoGxG92taOmeM+s/SecR7UpKhVSj421shywDpMR0+ZJ
iWswtV+vXVrIwwt9IeIHU64ugC78KtV+8+nMb7VaLWhzibo9ciRWg71TY4Gwh4u3PoNPTTcel/7F
kHkF+YA0su3eyt2Z6zEMt7ok4xKFjJnyAUm+7WRfVeN1reSikLzSYY9aQwTtuIaEIEz9IN/8wUhq
6s4DpKYUM5AluFCqCfI+qFONl0qDhbx4SCPO0Pug1iulg8YyDQNKB4z5333G6+PJ6iL0Vc52KDfY
DLR04z+mgtC7nBfI+pCuJFBuA69/JZBi3BqtyERooDZ/jvrPVxq5l54XIBEG8Yw6sjwoMTsmPauD
Va5/EvK7Pg/ddSa57Yq3+Uzb6FRYhUG4IYa8/FUnRc5C6vaIP1dvO4ZfuM2fW5l+9FeXut0b/vlb
4N5sa4A8P8oPY6/CPHzzhwY1eUaJDgb1FNrGrg+KRT945M4xDuDwh03JErD43OChOW0c/vvmhmpJ
zUMkLiMDqFohWTzCqMBWjDXVMlf4LY3oP8vOeUL0kzYNYXNqQLPmn5QWkH+WEA3D+6REYTfbOPin
WGwzlk1fk7NLy4jXSog+2eaOzrvxOqqOwFBHAiZ3bGQRHrEbZI5UJE5/YbnIcDURF5oRCtNO6acS
qT4j7r0WyQ4/0lYLPuLlX+Rg+1Q0t2SLrUsMx/LxWfKtRB5lmJNw1XJWYwifJ7u1K5pW/B/61NEG
HWF/YhISsPJLmKBrw7FPQqdhSzxYfXT6k/ytFmn9PsRMY9MIJxbAxuM/MBi5pftOCp232xUfsBI8
kPLxiH5CjkDDa3RE9VzkNCPHWtGhe5rAdzOS4DIpxTGVAOb2ouNWgffiB/mzlxHp44UGmleG+8EL
PdUG3j1nl9g37e5TfUzz0SPSOdCwYBMqS6vw4kh15BgcvEgKlNjAI6KKeed4nfefF4bW3ZXQAT16
muQ15aDtuPE49JNkSLbYSiJdMNo72GjcK1Nqz94bNs1rzJ5iR3DiHFPhc0crdPfUEyOO1BKaYig+
+oOfBKFBcj+ZiHoqP9CyViozrJ97HcWYRYioGwti0YFsirpp/w0O4nfPgffjh0/Rgec9RtvYA42f
Zf/yQuOhKW/+3G9zk5c91D0lW+TIvWPJk6rGOMa2flG30xOokE+IsfFH7I6t8sdtEiQU7j/t7dKX
SUJQAu3YayPy1VGosCFj30gyLvuX28bSs1Vm+kAPa7UTA2OkpXJ00ecdtaGgRTBhd3gnFDncqy9V
YPBslj/jdC2ZBLZYLtjknxNihbu90xVaQbPp8hcTXA0++1GB1cv9rpPSaqdzVmZr39/TiNiUo7Uf
fh52k3U7ic7lXyLwpqrqkUF9smWu4Xb27nbpZdcJMmj8UgvScCXiQ/WbmJbQee1NMrpcQnqKdKel
+aD9+d8qSyufDcPpRl1tRG3sPiQyyf+aFMLpc3v9iqhqN5wLp8vp0Fl4rf/fnUf1ryAGt/FRF8qR
4pMW+okmX5b6qwCgYDZAE5Rs2sZrlJGiZZW0yzwdgkvHoQ+6HdUms4zNnsLeRZY7QlLigCyJGtBU
mU3xB4paoHtfta9wLzoL0JS4UsVGRYZA5JKNXGCSPYa3/BhQPutRAojODXkLPEnRqzOepff78s4b
PlJOHWW6+qRb7Xb+5+6XU6UaoFaL2Ro8oe7AtziFoZf+A4dH16xjzJQYyCUjM3w82VR0FY2AawKF
rFQGZuNm6ajEGpI/h0iuXw+WvsiL5I4H8k3encVF7uDwvqF2VVznC3ynSKYf6+PVmDuVSgLwRac8
At3aSZyl8ItlQ205gLKAoWGM30wr27qhr3tD2nW9kpm3rExerE202m8p8velrMqymxsY8cWDpGck
V1hQxlJhjT/w323uHDi5KiBOhQ8q6/HvrIKu7R9E6ze+gUBBrg57oo4dj3RD/YI3ZYyq/MtICAnC
ANfgVSF/+Qc24IQVwSAzAbXqwteDicXwPGXeLs85v6ZiE6X+nwCpTwKlDm0heTILv+ij6oprCp0P
uQMr17Ccwsn3sYmkSQa2NTL+CZXGjxBFXQYj/esUPkjcpCIGmeH7jIKDQ7UlHIhJqBrC3Qp81NjA
WSBqKeeEn+TbinQtxmnIsXQtgcgCw5uphLGnWpgWs03W/Hcn2LL9S+5NdGGJFY8dVqRIbmpEigdR
wjKcqNkVRN780kZxLupo3tVs/dFJnCPhePZQwqB598E3VGdFuBhXV5sDIBaCXqoVe1QRHHs+nUbd
LF2vB6Cmh0pixkC8om2zfffcJEHmvcTfWgno/UazF+oUbWXT+ZUc11cEMBiMrRh39gn6eYcFs6TN
j6yma5G3mu771fE5eDxZRGZcZqWHIXQ7Uz2/uq7Vpt5yB0aiaZ7C4fAVKS+wODR+5fVwHFF4kKgl
jg1tukNyJtp3ddHakgilDUSfYGMgNuJaLvDjK5+ABx8i1wE0NW2YHVcx9Wwexy+Rv5eEx3xXT2bx
UEuKM/O5JlvOJ8Y2PBOqrtaN3bKsU+aU8T106KL0cG4GLSHqlqngj8IcVA4dTndxgvfC1ZgkuPPq
Ig0yC0KiN1HesY/NtZvzrb7C6S5iDwwGVwKz65WasPVFmsbAzYnhdZgfVG19k61JepdPElDuyc6Z
uikQAOJoXo9xv42UgorrUX1JU7AtAqzkmQdRddwjKF5+LCfzrdChjjqUw3ls+5muoEvzLu1xouH9
S5bDThlxCfH5qExFbcbv3qOc6+I/B7hInP2fU5tZqZISMk+3mfbn7379IajKPCLSvWttyVLl6ZpT
xCD6hoj+bbILhAE2FBBcI3RwOvK+U0rnk5HMO185pD+TpZnJBNnXFZFDMtrpxehef48+sZPLwPyX
AZkzgNG9ol0m1Go5SsKG4SSCLUwvChIxyGUNn3MPW7624sGbBdTvMuIfQon7bohcgfupiSw7fWmu
rjYsCibm8C4J93cORMP35LilUUweAlq6pDgUc3FnX/N+W6aF6Tz0/byQEqceF8423VeIAmUf4QPv
LiTIGXZkYRmP3d9HUmw7jYgsUcBRQWmxgkBpyOeVarukMV3MXG45Hj1jTB89BOGiW8TUeKSptQXW
3rfdLOiTIC/r+HsvULeDxdKXI2k+f/MuPOuTbaP0RcBtT+lWfSbPLUHZKk2rJzbgmsPlMcaalj0s
P6nr+7b0ojWx/XQ9YuupcFcEeuW0MuuSSMzv5hMzQgKiiRU2AnmdqB0RsS4Dw9ojLSJYKwGh4ZQC
N20SK+JrF0aZ8UOCuE19CMIvJIzct97fO0spElKfrmQkwBoYWuqMfGRtPjvio1g0PfxzYWKY2tIr
jGYK+h320MS5S3oRIUz2oGTYeRNlD0rkO2wSvuZnMk4HQCUpUGrQahfELL/u9NZK0lBaX8EMLKWY
wuxTiJ2EDZEcl2kdbGoPxqvo7WulpcymtAItnZgE8ON1eBWrLPlM4hYSWRbEL/QfxdEfKSVoP5cF
muHahUFkGpfgbo1Zp/HBb5zfI6ws6Kxwf/o45B6h1pxKPYA+ksxFohsfnhVZI8qHpUWAB6HsnooD
RkMpYj0LOKPkXZYxhiClubFO/lgOkmABkW0BMtslqH6xMgpGT4nL3pSsqe8Alo/udSJqcRKue5et
a96wM/gFmU8HdY6tPFhnRvahoMtWQtWOks9rkksmWODhm+r7/thPoIqgNtcHGefL/SOPEbdhTJKr
nLN6fU/TJtEwd5yelBjI6JsDqnY3Kz/0XTKEr8T3OeAjDRT7MdYesJbXutdBxIb7KlKTUjofgKl1
c7Id+JmZqm/mIShveBuUxst6wooSzNimdA9OOxW8+lraLI7vTpYdFwAvpI4X1FYjO78+CQ+Vlbh/
K0wWufYCn77O4Iv7Q2kf5cOerr+ZlCDrGZ1eWiyk567oJ6eh0J+BIHIs6GcT7NmrUxZvAoA+FBkZ
gErt3WXriCltQitDP7Y0iByXMbn8AvB+3g0CHPovIdiL+T/1FgPESrnUofvwrFiOv6v8LD6ABq+r
Ddq4sLBV7ptwQ9dHY4nqryO3PtrHlKUu3rFaKi/oM+NtzJIclTIf6+KJZvhmjfRso2pU1hBHpEXP
/l+rB0LBW4L5Rqv8rt+fqyVpJvIdloO4YcUMFq9+ZGRglsd02h4mUGZJLilJxpnHBPRCwkhtN+gU
l9RpEGmjIg1AQWT6SYqF3aoQtmyKQ7FYvEjKeUDlUJI1yMv24KlARIQBOM1sKlBdTs30AHkAum0C
XDVDBrSNrmyScH7Jym8JeynwRLKeycjVOPXW9c8zOLWxonqMXkO5YCPvx1D+Iri2AV+LpIgGkKMI
p7KVKJM9Y2LlD+krF2m7iOzyR23YzsYH5n6usymg7QZYQxzpfjbzXOP8TYw1GvWmrVMJc2CrOfwW
S/KS1dwK71j7v1xvXzVynpbg6339CAAPGqXA4x3gwOSum9Jir8QddWI0sG8l1w3CcDpzB/JjvfuN
cRDtFOn28GwZbsnouM7ac0DBsrnxTrheMJzH0J4nATIt5/KkClNfS7rCyIrwLy0xn4mA5gJwDT/K
9V4JqSyvuDNLKddIt2OHzBW7O9voO9q1E442VKj44iLxh6s9pESwwehiJdRF58ZCsrW862u1SupN
j979au7z6B6XQWPEoKuZzKYo7lrbKbgbhLImu+Jx3EtYpG1NbQGQrmAKZRHuOGxONe0swXztsBw8
wWGwmIseZw9gqsUiLipGsQi2t3p7YFb/tuqYrphW2qCqYXg5P6UP8Nvqhpv+sX9QvPBGZ3MwKwfo
iyj0xk1YALzCBCIV4eAzfJTnBArqUoeAKtDkmcLRaR4PpQzEPaSz9YEaL+80ITtIlg/bnPtjvxwP
DA9rjnjHlVCkQbCpbodR4YBfdG8nAS30HwH7hqwpIqErZbgXqxrCuKE2TRNXQlr0LSTqdZmsK532
ZmFn/MfcA54dwkprdHylzb8ELlGdrYJfK0A/dzT8Lg8kuv6Dqoctsh8VTrsPczdZPpb+yU2YnL06
rwRJD4tdojJUlf3wix7rce5pqZ5RXpBL3/qTYXktcgUmEbWLbv3niVBbR4M1ZANBMf4XotUQKIvB
BPbAlOCi+zJaWBfG8nn+mmwc89BFXvyDNVK0eLxHr5KWhUp56jtHEqtYpOJGyXTPIN1EfRr3nP08
7lphJp+AiMZ/vqIptuDVEVid5syZhw9+PiM61328Ed4f1B0S3X4JBRJWt9G63ztpoWC/dWK6Qwiy
M0la9lVLY5rILdYz6pqLejtlpGbCeoAwTFD3EHHZLuGgOlOqtDumv1Jrkdgf/9YmMISJAKuFsz31
9MGypf/80DdHSy75Wsg09HxYM945SPkjjmRa7SvKkbB6rHaKIJ4Naitonb+8qmlI41DZMS2sd7Kn
Hk0fWKQxTtPbKwouMZsP8DJlC8dCp0OJ9h3QWqnmtXBwQ96iuef1ahkKV5kOajPirf6Mnfmvho/y
Xi5pBgDZXqAO+6KU5et5qIlRJ31u+J7blQbnkCw1UncvOsOOV5tJSPxg0CCcJJB8YaMsp71cnGgY
96Ymq/O+wO68A2USlyjM+VXm6EmrUNwVcszIQhS/UKijjvSdehe69oiz3mn5KHb5+71JQ1PiaTVS
IM5g8dYuNiWJbbk2weHKV3Hbb2p8TbDtdzl/F2+Ux9hAiRNiTGqIKehmvesmZENqvLYbnKsYut5K
AU31WL4nSqw4YIynFqUCMVekT79V8H5SwMFxqKgtjiyFUkbBmpSSDfdSr2atDM0AlYHi5d6mnxSn
D99Lx2hxsZzcX9BjpVwrvJDe8WP5amYPL+GcPDaFlgVESevZNyw7cIbHe3dlcwH3Q1jVLErBn0DI
sgzfocbnMv4u3+I8VTAs+3PCBOLGZs0d0RxwIgjtWvxbt2Z6wVYSBXzaY4CHm3uyUTq3vXc6hagJ
UYDQsjwypeI+gDHI0Qzmj7gu4pmKCqPg6aEelPq8YU4Q/17FC/onWb8UH7I0WrCToXDwF51JYSil
zmgfe+Poual5HfieI/apz94I6c2d1dRfsHr6bbw3CjVmnMZ8OQeUQ4b9JcI9qHIoL7a/mMh/U98R
xmWz2Gkk7KmFFVdx8DxHFN473i1gGtaeyWAvMrMrpJ7XkWeau8pD1rrXQJv/i6Jwab1+Z4+zrVWQ
twRDJw9NAK1SEMBMxxfE6USiD7uG89QkDuzJAFZzSytdsVIIeBwmGQ6QbZvZowHFA9GYR5oGFr9A
2qdeZmGrB3Dwk24npp2VqA2FIMgfdIyj27Jgt4Dzum4HnY7FzM7yV3t/+JObgV1C84j8CDV+9FDx
kLu9d64Y+sjbIQ6aofk/E3uEOa8qKuEhY6lL9NnAjRD6X1Z++54rDmIAa9tEVGvi5EAUFwIoln1t
B6bUPFoegkzKZ4txrAWR+X7VoeGyJCN0hgn5V+kW2PlKJ1CBMQnsliaZY8UMzZiVsyR6xHzoK+xZ
uACPN1iUk/4Q/KVMcd5VFUq3zrF/u5ZLzDqDlfIUFS0L9AT8J6sgOjTidvdzC6ninFsDhDw/Yas0
5ihBCYM+8AnorPApJ6IRKl9/fF+TaZl5Qg7xdnGKq1ik/2fLMrrO/CAv0Qz+tfgMcss9ihW5VtAx
TWms/qCkuyURJSYyMiT1UCpDaC9caBB1eZSF0TJJKyiqfYRXZP9y2cF3WUaZsAjSqX/EKJPCvCPu
FyadaPohIieK+wFZieqOAmwI6537C7sIiGh9Mxb0++k01XBu10HWmHTZEIMcajoN6ooAqyAwfBus
dnKMzcvGLeHvzOoQkopv3FTDGZByIx3+m47sgRfE+wi3njz2Y9C/QHzT29ie0rQMCI8fJqKJdFIY
2P2MXnFYboO7nJE4alNNz2VVDpIBUcHamkIv1KE61yknZsW1m/Acc2+kYfaXoJ1TKZVabsOqwonw
JdEF/NzgKfQRFWg5BBAEiZlVEpBUvFmYMdBGGmFQodU7juIGUpMvPV1E8oP7v6dRlxmYu96rbl+O
EwvHfJ9A1yzI/3m5aFPzk1l2xV/onu1ezZk34dk3mEKr6OMBRXxNIhJQY1VF5asI6b5+/JsTZ1iw
MdDcagOFUjM4e/EuJJ78cYBbnlD817kYboCouD92fXuOZgQbrGyUXi5x7gDIsftb/UvI0PYVanPI
ZSFFdBtaHctIYt68CQfC7sUOUcYf/B8ZaElaFAKwD3N8aJOjCAXDJGN4GYEYU/4nyHgNxFWaoV9N
KLSBcb5c+xoXaMuBS776m3r/sdWVc2Cns0K27VBGZKxltD4OXvVr/a8YilUopB9+uCWDoMqNXHpb
b4hir6o5PDi+S3+/GvlZqcFSky52eSsL1RESH+aHl6UtBnV0ZT+iogp83DF8B7EGdekTuOvlT8vH
50S2Un4cFdW+SxuYcOGvdsGYqGnCkvCcaJJz2OgZf75rvXvJvvhzrnEJhwbPsZd8hMbrtD7vRNLR
Lp0p4PWs4nfYK0MWFELIMLUxhcrvxq6qfI7OmNq7Zzs5pFLf1dTdpnYa0AZVb1CXKYwtuyKDrOc8
efVTbxEk9jNbEvEwtptAzPEV/OFrr1VDJxZIyxvvfBJjjaa9ll2Bo0o/mLP15SYEemVnrOdzjWE7
Va+eM3p7D9BQmAaRcNS+wasn0nBS5MRnrqGr1TFX9pJn92AZg5p+2LT09lFIs5u1R2xGX2NJUvah
aW65QVAmRO3yBMAVS5c0geYemdA7tda2cQejJgZ+GcwGo9AezloqBZPaKAr7DkLgzTMO4TCEMuLK
6BrbrmRyQEqkza5uaexheQCQ/Ky5Mzn8/aiVtrbTOWNyplihG2b+ng3n0SRukRZG+bRP7IdTNWzr
WrHkrHN+1qD26yZrFhIq6fEKAju/fyXjARWcYKUdHu7xPK4PPsaSH0mKUoFNtVMJac5axqUXy/z7
fwJpaTqxJCGKVeyBKX3gZQoDYTflZLkdSIVWgOi5DfWwk9x3VFf/RJE2HuNxPVzCfSvZsoxVbVo3
9AiTicCvtzVx2fgyMz8YlBKCXCs5wirnIJr46BMIxQF+ayn/B0aKuTmmC3l22oNEr4BnTrsEt0/H
nZ5PvA7fvYknS0zaERg8uyjAXtrqXe7bHJhI+cfa5fD6bKTG25fAaqr/oWVMCkWM2oHA+YThLqm4
s3oluGZ4RNGSjBcljFzfdGK6glAxAWuo7oTTvtq/OibA6/gxu2USuciMNobUbJ833E9thcaJ1kTI
/+YQqL76tL3+okfjkoP0woPHoHV3wceVuxU/UD3k16q9kPwiyqJum5y/rQkO48UFl9tVn950kQzf
6yQB7ypBgmg/16rtJDWIhQ585gYKhFiDKbuJxQ0Cpj80+ER96BzOCtvhdST7DsNDj3gTCyUq4D55
9kOBd8VNu3e08yIFNRAfdilv363raMWrOqimeXW8cfWhTJhdDEhAXVx5XHJ0iwB2l/hrvJU8khAR
SpkAX96XsDzWp8awxmqlEdRU87MhRSa/NEP00shVbc90K5DsvkUTPL9OBB6egoxfYc0X09Ld9bVg
l9ExsIG81doCby4ae4XsetF+T5p+oMSCnIX32Ut4I+/MeCq8EphpOmVVQ2Fqnjzv0rcUIrR97LOU
doz1kmwX7tK4ZXtizj6EJvrqMQX8jnS7cvTrjqUUwb6YoXgJh89ojAbVWOdyWNjdHP9VuAVxhq6P
7oUKthNhtIZyN9+ddYXwjNPnu6K2wq/iSWdxrB5WS0+zXgfEqQ+tkhCjIEbtnGM94Au3+0wB/3lv
ef4nTsgQPjnaS6d50qj4Asb27KG/1xecmbdBGKZhNGIfRO1R4nkOCA9f5yWOLzQUYFlhdYVbPNbN
NlzeVWnnXkGQiVgKsXNsCzDOEDiJlNRCAJipqdyJmXv2T810WYJY6eojd92WWPVRj9+9GdhRPZt+
cB6Nab0i355TyAK0DqLYsYw9sk5F94ZeNMSzKqNHtvEROJGqAU5t3+yDX7icLkXNI4Mf+oMUDZUU
+nKakUvCyx5XQNI0yaV5RNBexocaVCTKxqB/uEF6OzSqKfsRglw2Sxsg+RTuH8a9mQk66vAzhene
vY63aMfJ21zwvipWgGt4FVuP8V2ZCPvz0QtHxLILIuETvcEDc/kZkG6DLbkbv9A+R2t6durE6v09
pMrXAdcExb5rWEMUq78Z63cXzk7PLf6zNJ2f/A7daL7zKq8I0tiQ5NsKNWtfuxYTO6EfXHVf+Djo
d2tZ11ZikQC/h1VEPlJIG0YcqcEcqrrRIx1iFSktB2G3JzL7ilWJbzUVemNuLx3A3ZNEnoO0NgGT
gtrBW4x6Lv4Zsuw7hNtC4W8P2fxxiFPzDtQwmAAf4hWdmcxv0ms5dveISsbe/YofBHZpB+P3kbrH
m/8FymSPxXGAlgs8UPwFUe9UkTPI52JGq1S2zUVWR8jEql2IUqcxsTFJDV+VpGChU6Kh+MO9Di0S
48PDygCZ6pXq/GGe1ejJy3MacbGqboTQ7u4LQ0xUFoNXAyR9EkGDzspmauVDezIfBCQbOlsaBidG
OoLNaKoj13Vz91Sdx3IK7nt488jD7C8Iuc18aNchCxqZZC8sNLh9B9xfoIbrfbD+6LQvLkUK7iGj
F4roi5dK1qKbOTeO3H8M60LssMqRbaKGDOWCXWjmgR64fE5GO1svyI4HAsESZkw63pOgeoYafw6v
IWE6ms6/MWI+55GP4VJDKQHLGQSI0xJad/8UsjAhQILXiXK9b03aLExkqmre+h9bLmJTHwxKWoTp
G3oQwSOZN0OCV49woJf8ATHJ1gZreBSxW9Xu5GswjjlW6EDiP+QN1gGqFzAFp4qeD2sYIAYK/lN/
b87G6CGfnumhIqxtkuIjqVWEX1K3anlpZ8rEmh1AAFJcXFRxalblyq0+f7/KynOANMdf+bZaOiRN
GhXmqATnaI3aVYy6jqjnJs9bB2XU1delahYVjuoyIse8xfhmqCIy6QM5OLDlEgSzVT+1UPbB8BSF
AsIdaIGUOGPymkWQHuaz+GxNEVNjZEKUdA5XZS0CqKLIiu9Hn7z7asW097ei0TbV5pcGguxZ052q
FND3bUWERV+FHNHNF2mN/1wV8Zl1a31PivW/Krr+c2SZbArq4a3ych1oqEeWrtVInYa2jaBFko/N
ISe4AsJULWgP2Ao5zdCqKHIBVeDO2jFnOIFb0pW3/cXnhA8c+CqAPxwDRo4F5bomwduLr5hlQMlz
FIYnGrINwJEvlmHG78pFF57uH9BwwQaH9T6cK6ghyoP2nZ5xnV46V4BT5oAvbWVgnZIP4YWKQ9wA
0OcQ7eQKWl890SVZHAoA5vhwOyD1OkLgws56ioRKGX830EOp4ztRbLAgn9rf6ewkrP9fdcGopvLC
YJl0kNTLzsON0ggghl1arkvIeKFJv9Lazaw1zkOXlLfUYVc4PDg24Ri+/uv2hqxNCJVjcFqmFPEY
3pmVv+mGbwYJWBDlAv4ES6PJNWITW4TtVMeTRFgjWXPnS6xWUh0eaxgLqRHDx/Rlrj0vAaxxvX9n
kVwvt2LK40YBFQxHjHYU+wnCKjCXyETlFOpVCeBD3IqutF6G1ESNno8uF85/XuPRjkHUM8ziVP7w
RL2WhGJlCPAHidiOQgwYxIy7Sc3L5E0COmOlVlHEwS5BDjyJEAvWkKEY7HTkhMTwuZmI1IgOYzmz
GDvtq1Qc4q/4kw5osqm+YFh4lXnZP0asoahk7wQaB89enIOKLAqySwmordcyofH8UL053ydeszts
UiO2gmrDNEltZoPRcWlubkLfjP2FZPPiZc0TR6YU0uNzVR/+/R0lP6elwCy2S1pV++NiOiYTzi0+
4i9KggBxydbn6MwGy1isJzm7aIsPMhb8Hw7/KxkgCyRICT0RoaGUTp4YH6fyGxMyAPdSHvis7i+4
1+kM80mCH0eGYfWdCEEFbgBrsYfSuCH7w8atHhIx1OtAfkBj+r0Y16U0hC6RLeti/lH23toSEMgK
dwt4USynY/qqmWqgf5cJ1y3ZXxTyDrojWfGO3UlesGqrgrUzvI3YVOMRaX1fN90IEFeynbfKvQKd
Spmbn2KCyAzLOeNfNwgKqWEKEvo3zW7GxYUMasUEOFqhfD9GWoBHMHdWd0Ba16NNEBykcjv3mrQP
5ViScluvZ+AJcw3exAu5mNihdgl5t7KnInwsrrx54VOWj8HGEb5pxud+P4yR7CBpqWEGpj0yjuFS
5O9g5ZXfLn6zVWt91aaLkV+nW4NsKwhFpPpD3CYF33PGOypTXxw91GRUAuwz2opN+7n37E1OFgbJ
LaYlMa7PKCHJ44G3hQrwDqiyCX9t77yqYNCs0akIJz1zmSCCxx/53LPkKkNropdoqakji8lioj8T
nk9jlsKMX8pXRRq+EyfXBgRegcr7lF9r8MIatNTrmdWN2eWyJQBLYo6ck+xYf33T8xuCxXeq+ENM
RZe5p/gJtc8dckBNJDuKv7RKicfrPBupZP0Gd+kzxkm6RPlE/TaLhT1FmGRp9dbaDm7kwsqEwb2s
v2K5FxLXHHfTuyqqB6xmPdzv4exsLtSeZNnbps4cu+n6Mf8LdmzORwTpiTLFkwog/B4JnmZhP5/X
848t5XLqbgqnGBX2TrSrai5qdoS88Vejf/FwtkF+awrAUWPEfRfLPPnSIqalZCPAobJOQERRgqjV
6fNiqzxg5yF8lH3QgklgyC6ofarrLc1a+bbPZop2hZU9GFtt3OubmvwmovKqWx75BvEorJOUxloH
nosur585itLxsaNFPLD0dnnWropY8mrBIBhnq0wvkyaaA0qcBwMMTXb5hjdRNSldzHIdwTq9deJU
Ri7MTP+gyyqcng3cTHFo0HjBe7NumJ047wjQdWUtQ/FiyNDWakn+e8L5zrYFbt1XPzfawT7Z/s9T
Ny3NuNspcpG4IAfyujij/Ll9Low2tk7noegZ/7hdRcf3UU7mfI79/kyvCHkF99IJD1W3MSI/15/i
0DkkHkIT8U4oKmp8B2VIDURzYWC6D88xdvjtwIxMs7yEm4PUNeLYqJsJxesJzEsXkRieGmnj9EuG
bM3AJNlRULpj/zuSmNp11iJAD3+oa2C5X9MakkhSObjDPrGWeB+lYdlWUwx5flTyLfy9XKXkH/uT
calRpuAh0JTtzvENZn4AHj9jUOCf9rpbmCjpSz4vHGB1UOVwXIQsTy7dX5+xUxrKhU1h8HEKReW7
B/LvvsObjaw+uKlKEJQH7fHnG25Z7Gk/0WdKgHxKdrcV/R43FX/LHT8IAtUdCrLlsruvX6zK8j7a
rKA1mP3LPrN3udHfZi6IDR3DqQzp/VTInnVaXNrVJ2Uog2GkKsKVRnUJmhRy+VIwrPZs0uvN8Y8T
P2W5RG62Bqlpjld6/TenfdPOISTNKpnHoVjyfDBVfiUNmC4Kvsu4jl0J8KF8r0mbcpschTudyBlX
Y5AgZEzaGiEebpZhFtvaRWK5pSTXxv00jQdZ52GRVIJ6WakyIvYEsLfu2Ch0YOIvgKdYl5SS88KK
kqzgLTKw8oqlVnofgfoZ7LW6RunVLk70LpGvyHe79CktX6Vz7hwni5vpg3s+zaMxhXJKV1Cg2crJ
ceshVYJS81BQqpp8zIrCytqnTE80Fi5OlMJge2w96Gei3ExBM6EaQK6DMiPnVPQrIaClHShb1hTI
pog1ANVHwCgjZYRVnEZi3dDuV258hdzyh1bXaCNzpuBb0nXnOaFOkTZX+qm5F/lNcXIPwUAz8D9a
Kdw7VVcVgVeAi4XUqM2wn6Zw1v7+X7vrSGl6qYO4aWQvafiAjuhtFyHRI+BlqxuVGakwHL/mCoZZ
/HiMTO9FT32JkdWczqV2ZKY7Ss4vhxsslAPk5wVWna2SdSXAbV1s0s2+OnsVGahV3t38vRRxVyiq
GGFZRxJxzdbH6GL631UzHYorWfd686xPVa+ibXRLMcL3Yw86VYoKE9eHdrDQ0UX/VBotPssBsKSe
7iYVtsLBqp++1Dnx8qYtbOoaeFKNhwztOjLgI1XcLgwXvO2x0fZV84owxH/tyKN8RJWn+czwlEdV
lGtvN6bt2pZ/zNOPvW5J0szowtHBApsz47nk2P/1Fb38ZiNC75uipl+wOv81AsFhnP2p8oLzOAAJ
JKjt55KFiChOIewtpghuYM4h8PBAdUxHr7UiROq1dVS9C+sn+u8PqyDzMk9AWArO8esY//XhTIHP
8nznNCuOTN/5d+APk6O0aKaYY2uGiWugrOnN4ksQLTrb1ovzVWJumBTThvUfbUBiqQyoVG3y8Qmr
ta1TuCNMaS/fbilprmzKPBhCgmlDy9L55WsMUed3+K/LnRKgjVaegTb2hp483MbCYX8zHV65LEu5
3i2AdeN9gUILijRPeTujrKDrfCRQThE5QuR40886bx37SqN+ERC8P+58ebzVTN+HRsTVTWg+wQOj
1NI2l1vhDxinmkxYvcOei5WYkWUiWZRbcWgFyHIvo5ihjAxHMMP+8m50YzG7hH1YDpiYRsiPpA7C
v9Hdl1SHRjp8tIrhCwgfdZdR9sq8cwIB88F0jSqgwwgz400FZATcqnZ98nVXci0ad1YhGFIdXYBc
j2lBIdxTjzPpQDKT+gKZQk0zyzefPyLztQU8V9wlaObBH1eGV/18todjq8JcYHTBnB9PKrw3DOln
JVCsXDylNpUfp4J3IWI1fEbZ6deWZULmfRezUapvyb+0KSo7OsF71YAmHVOBkef0N/TdH+s09Nn+
MZcLe0lc5AR3ZTDgzTtE7NYhVI8DMnj4z3D/WExrMhfiDqTNdra4vMB7KoC8TQH1GlTTUxcJeR10
qob0rW6iA4xv2p3sOCzydb1ke/eWaui41jhe1F+C6w/Ylh7bhUL9Z9iYpJoPAzXgEpMYlWp5/t2y
jwsUtIkY6JCCeO8u+7CPh0Wc4Q2zFe3C5J0DNmb4BUDpe2St3DtWFXpk6ZZRKNUmlr6dAyI7dn6y
PwB7D/8AgA8BNwsNEzH8VB0o+3Atfl058W+xFoHwbht77thGppw46uaEEqHO3ZDBKuEtep3JHIPN
UGZ8r4Oc9niYFIwdj+UyixrqncD9mSFdr1L+xEOTSLZpBmgqMgN6t9Yl1JXlo3AaMPxUUQgDsEev
y9giB2M8BxEbndYQ5pTAe8/QCdrIzxGO8NXJrW8pfiyfccftpZ47mpLkXz4Da2qUoYK6J9iW2/bX
cwec7Ha6FdbkhrUb36owRaNMxTp2Ip4apsX46FXIHxN+fV22sH1/PRkTgyQu7xUlvZfz4XSR40f9
Q2F99msgo2OERpiMORIJ8QyzyjZoOKGycYI7uV8++gwu0DLAdiJt1GupiMcV+PfkZAv/HgXIIagl
0Qx9DDr1tZX5/c/i/y29d1o1002hLm22UYgcV7OGakFuehYFW0U+AHCTN2N4/OSZ3rMcjLZFZ5JO
YEX4m7O1eVrkovBZoUxTrIuI+iUdOt4/rqMhMZE7bvx8QWb4ChShmehuMxAmGskP/g1UVLFhxNzq
UCsIQ4df/lgy7Y8uW8JbGtj5gcznnEJck4BoXeUnCx7+V8tsn9mVDZD6qLw0F5D46Nrrb3B+nUKU
xO7A4SkwoQJlPWG+BonMloMKv6RpOGoaG0jhPoifZXXYIBrmWEJN2xoe8zpPDkAa5Bj5YG6wwcAS
mWPNpk7RKdCrT1en+qSZ4jTk4iuQGQ77hSSYBjGCSR6cgZMlN35NlO7VqEsAXhWc+u4ylLxHxcci
ZXhbPq9dPSpQxHB44fj7jCEm+K93qR3XJraAbCGfu1XkbuugPTlHzjaFU7smcaQ4mHpGCCWiaKNt
orQ1KtnLLWgthfAqj00WWnyO/42bgQEWpfF/sMqSVxxntOxt5iCVmax75aVPWsaHPzftTyM8FvPj
49sq4OBljxxqLkjJL/jfC/aYXdp/pOXc93kYpmp1zIQYD5HaC9sjNdvZkRnd/Mor2H7VFvmIVg+u
wUCssgA4eaYTr0dTgeFtDgww85DTeu/B2237uol5zfUm9y/gsvjNF1ijRb1Gd/GjJjSPL4gu6rQ8
vXtsQuu32t1TqPlxuXpr9iTi+PnOaDdsJTWIYSak1uOCYgOnhs/QexTnKrF7Htktwm7ldfQcJ8sa
PWPvM8M4CwBGheNj9sJ8ykwkOYfeeUBCwN+RgmSeVZFBkA2hJPnLlOTqJcU+oUA9qtMzBfLLDdmn
xzWN+E82DTdJA5lPQ5UX3WWg0zlhMW2fIglBBc3+/zCAIcRk+1Dtf2HdGC7pyWKa6P1tWaJVYlid
JAJjQK+zqgJUTplDla/RSY4Ug41GOQ9rWJQs/G1E8qiSQX4nrH/bxcXEko4mYRDIxGx2uORgKfJY
lSjz2/FyAf+VrLTwZSU2uLFPBmHK5OOs8fG/E7/wzzrGayMedVfaa1Z84L5UdD9DjwbSHG6GL4VX
aQJPxLM4AIbkmZqqJm/CWKhhcw6HcqR3a0vk9koFcqtGKWc/yBKNs2Qne1PgHXqaRDduRfJw25sj
g7f5kEN3AEd+Iv2pKJ6HYxXJkFdGdy90P3SWB2EaJShlZT7N9lT+k9NJcnyRVxTO4DCdFBnFXnoa
HwFVoylk1eV9Vk/fuKm2OdBqu4W+YK7GCJJxHh2TVzrRIHNEXHJNjMJQdx0xIjfa4S4vjH9u4/qF
qeZBD86UUMNu0VhnY0gSeQ1oTucm5cSLQRx+79MDnyUBEmL2by6c/hKjWCCcJFlQ5vRx/BurQKdp
0j61c9TW1Lnw89PF/AatXNEuaqYVRev/HiszLPZ7pwycscmnBQ8hMvXfS+MTvDwLej9AInI8Setn
mnArYqUtzU3HYor2TauNcZS/eSAczUVqTGnwyFHWBjQ/kPHlkHzEshCNjJzasjfNYIETlz4sZG7L
0ftnuxqCeGB728GOj81LgFCQgGacE6Cvp0uJBz2odCagKRHqIa33GfT6QxRcp46W/8Nr0bvT+xLO
z3RN0/jhXA8Jsc1CH13L7UUyAYN/5UaX9bwxu305/wGNVaVVCh8r7sgBN4k3W9n7Q8Qs2hGoneEL
kTaRsMxlUrJVmRDQQW2u8Md+NLfXEDOxpuHEmA7EVYQA5f5d8C0WTkoO02PJ+LrKH3dWGuaghf7X
LWoCAVxWO7ghGXmmgJ/1afZeEW01qPJTn4c64HF/UUB8y7HUxVqJ2EbPEgLqboQugn8PZuJBMMJY
iwN+T5iMgBAdYzMJqlTrJNj0cAAmuBHHZrqOYYc+WBqLsmbcsogV60UYDi3Ad0uxI5rlpEYziM9c
wnGf3kI1EYkqkT255OrDmL8heqZf6jJfMB9EzOURZ99JmMN4srwkOvP+K6dJj9OZ77yeQYcXqqKR
EixM/YunDN2KEmjS52hKtH9cMRCHuUnv9yEuGLUi3krBD3tyFs31Hxf8fvJ68TNzXu0aCn6tzsM3
oQyW5QcZmFlHYtGM7vf3YuPWBxYagtDb/StrbUN1R+s+ouoimdFiQQzbbElgbydf2t4QvgGGTmXt
buBLd+jKpay7MKC2T+uJ1Ex90GlyjuOOzi8Kr9UZsMJRCX0ur1S7yyYCO+uQlTsPqLOa8zPKWZN1
t2GRVXtHDEcRbOISNLIWja4qxqKaUODAiU075E7R0GuFyF/ZtnYUBbVq+JSfVWeBpN5dApqAMa3/
irSc4ETiknRuLhYy9hEFEN0g5lloImNRPubeBza2Ct6aKX/zUkHntzIGwDnkyka/EjIiq0GraqCD
GSCvKbw+oYGfn9Wy0it2ftA7MOwcHJUDlSqUqmo0oy6JGn1SXp9CazRujKyObN80RYgR5fgbS1f6
FyPG4NbmuDIUXv2DCpX4x5RFhDNXHaSarrst0VUotGAskuslQOWsucfgJzIauH+CnQVn7Zrl8861
lDEJggujnq+5RbDVmyx3EbtzFneAGpw5HKjsk6IbQ3/kJrqqArtrDToa0n4YuLNeicRfJANds/Th
WYB1MFF7H7H0aRCQJQy8+ZnKSx+Cm+0wR2nII46tFKYMMz5p+4y9uBZ3UQ2cWu8nmvFba/vrSO8v
rBbK6JrP1VWZnVc5/63Uj5EcIp5VgtFAHTLm3TguzxefSEtxvyroZCPCh7+euD2/XyxYmlmprofG
ZSiaFB0V+Lg8UoiBN/8VjN/5SAeDsr/U+nIjJT5+YJYTw60BhmqZLLZ49giPq8usZMugFZVp59fv
tW8PB0ztFCZQDY+Mqy5XXM00ESumSZvLuaz2GjOif+BWsgoYMbhS7EvynSxp+JjWEmhCRA/Eopel
K1qrnVp8D19MDaQr0CBr8g592KOH9bMQ3kdLEWOPyAlKaPTLGhC9BdlNp6dHvma2sKj76+3QkWwX
fhyHScM8+tJUS4y1/FaCgFXGmaHfTT758rEEYFrd6htJuxyiLQFY16MC5xbT8mWI/OoNjnKsTa/9
u+YKPpx3kODgCR+Sruo+TX8jmZVyux+4Cx9cTZOY8vgSgejV5yc6S0TsacUkOEMaXUxKqYdltK4I
xNbqbpYDuCrURljUHNCk8eiODzDyw96WLv3vTuLSFr7b0emls6abxiAC06ojiw/HrWwIRZBTWXWd
dhzBl8YifHsywjpG3qS3wJ+TOK4HPDCuzk/yln6zwqMDeFrzwfQpBGh4e9TK1GjNbN34hTIQhOdL
CzrTm3xgQfcsTlFb6lLGM/8v40eFnZZu9C/vdS5nGcuY4H8Z5b9fGoG3xbttafxhPHa9HwWr04J7
S6BCSLeJNxS58wGc5jV1fzBPP0DOy6/V3WEoCBOyI8YnTORLKtMhQZ9PXYDCPtqjzs81Qra+DFwO
UnltiB9bC5Ee+cLAIzR7Lu0lCDlEPMYA7kmHW5mRfn5IjykNGw2qC25zCTildOROFwUUcIT/HOty
syrr2oOoZAgal2toXzSudPAqqq7gTBNFEsvtQpdZ6UHfhwh63fRqxXLF+agl2M7l778EuayPWGrk
po9l/4WSQir/tM0p+429mb4nqc28CunVmBUevxEjJdeGFTnyldhGG1xQCr/zuG4Dgn8nOPX2f6+/
uWBAasqQwohIQSQLEmItTX38AkSXf/Al83R9S6MjHfY60aqG2BxFtUFN7VCL2sQdRIjdwZsjudpE
XDQE65KYeZjoDjutD8pEEfG8v2QPOxermX7mHJzYgqARGoiQLIEpWhM0pbi3RNM6RzQDIq87si+T
PSCYMNIThjtwTDd7Izcb6aMX88c00/VAMJXLVy3PVEl+EQKyS69DRK20bU3jqKBUJvLT+AZ94Wiv
XLMWHeVrEcPw/U8v633DukEw+sno5LxLNBsEnF9I8MPTilOHKwpMoE9MacOcM6485RlYfhbHMhmo
CIUR4Qd5gQBktyexPBUa9Z+dBigaSlcFGnEpO9UyEWqOecDlLo3om0fowbq5GpqmHLdn9usCHgHU
s5PFYnSGd+JD5cpM3Y8e20WQlVnYPUPFyQcoeRY7ZN+GBxN3sZYf6HS+9PSiDQd8NdM+2g/jgO+o
fO7Cf4r/v9sGm9kNOciyzG6ONfhsFB4vkOQKBOTFMvOprDmw9uqfrLaUmMP3woAk2b0A12WjC0OR
jDi9xSMmgWCBeVw/3YgVSgGHfLXfc/DTTa44X12Z3r+9LRuoMZhS6uFnFOZIPf0S4x5jmsIZUszO
e4p3+ryy1ks9ucwYt7XAnKjC1fkZCAJUx205eVGkz7IdxsEptkOxLrk6dKaENzNZn+YhDHrgxl61
3sM1WN+5a8hAJeHVTfRl96XqGwlGHSDSaQEOZtvnh1RwUnTmfAPU9NIp5rD/Iv9CIbddT76bKevP
RTe+jxcsLPmuGyAu7VpjmWnToLaxcHPU2sbtncS93LNk+8hWETy78Yh+RJlo1VMrcRj8Qa5fZq5U
s5jF8q1z3GtssLp/9xNMsB63cVksiTy/J1nsjmzmzIdwqRjLKjFgjGcNtUVg1kl9Ha0dkMQAUbCm
2kC+U/pOlLrh982Zr4z/uo+Hl/BfopO56ONZYKFW9kMZ071XVR70/sIsFxIJcDZpXFJfu2dKGWXK
TIReMYbkKeS54cv+wQ+EVszvA4vSrElgBQwlEwZhmBiuOXcZzOES+7q0c7VmV2EbQA5GbLUQib4O
uK595XYNWbGsFBKz1Dv/0mGoA0nqNL0WXH4kvNNjeav0Aam2nHFwS7v/WN3z/fOEdvNVP9IzElZq
LJEWkUBpBVXt4L4meJozHDSWATTHfIHQxfT9zleTjl7VAEgB4pzhPu5zVCaCgaAfWscTwXXNG6pe
2u1kXygXeh4O78tkO+JEl4vQOtOxzAvxuT0cvZsTc77tXG611Lajo8KzhVHQhzMtoSDTuaIAehNs
h5Sn2qqwya75DKVecgRkiZcT8fVTzQuc9KaW4PYrJdpqLwAO3e/BlLyz0fhEoQgFcMtaPw10mH4d
zszvhp43n4Dx+56pKrlaBNoAfo/1zUwvkYyYl0x7MOnGmoH6pTqZa+MeOx7sCaee6UfiKHE+b8lx
XhuCoNvg+dt8aTF5x2caGQjLh0WtKwACW3eC42MmZodDQD17Ur7yfAIfovqJy3wEJ0NInQZ7VZ1Z
oYozsikBHpXjcYPvPA+QldjzjHpZvjR3aiuGr4csvpJLKPAEemmwo7j3wU5/1UdxtAVAz9Z9f6zc
yF/qNx36W1elU9o2ePIhXOUqZYCbKCWszkiRcld6ORkioXjDSdmewPCH3Ghw0DRCF1Oj1HfMBj/Q
e1aJgTm1fHdjc2JnxSqpd+PWq67jeZ3n5m+MrIYdNpTwaJ2zFwRzkFScXmUnJI6lauIR9VbU0MTt
kyBTMSmNWUvUotTftMwIpps/NlRxG65X0mJ/KR5eGJxdCuV8Nuce2Y/8dfL9TgnOmLA6OnbbYRhm
lShYTyoF+fZcAQ1pmNgmqjw9GGd/Ogy8pPZ8MenqP9guj9QAiFBFl4mLZQNBBUo6L3nwRNtMugZ1
2EneExvMyJmTH2eodHy5ltxVbEvzLf1+RQ49XllWKbka8GJOd6de0jkWV2ntK1SWz6o4dXWT5NUK
OaOLdY39UY42sOeKx25UxvqdzDj/xSCbUSO4l8no4qangbxeGHLPfoNPGDO4PdCNlI4gu1CQiQ8n
n/e86jxRf4D8QmAgb2KSBKiyGvumLdwq8RJBKH5mwBRTrZJhjNUH5tx60U3PQDTVL/FtzvsQXiYc
r+axrf22+3xZoXI3KxTLFmVV6GM7tcCcX/BLVrlv8XuYDan4MKSzqVSS509zdgaqQBmowJPNdIU0
MIb21+nBUuj2RPW02KK8M6BDjVyWpY73Gy2xIQPPhZT5butvcvr+VPpPtiZAoeURwZ6lxQihi5NU
II2QVW4C7EM/Vv+WsfCeHV3SZRSJ5Rm2BtNhJ8XuZifRKgJ4Tuc17C3w751mbotzkSzU5uQ92eR5
2WE2j1mg1iZtwUknz6HgUYEi8/yKBb8tleY0t3LS60F1nc4kGERnV/T7DakmiCdb+NOs7NgUcjtT
wNmnxXQRyPIqVAJamu/8erS3vlpp+wJ/aPbEcfxNiGM8tpTLNYYoVTsUTr7GM8c8O70SABu0bhel
jmDE3IXW0aGvsOVWvBWiyB09E8l+VaN3UFzq6YxLqj5P1gfB+c6dTOuuIsDUKYrDrndID7bQr0le
gm9+mbZk0p+1doqMvNHd0Qg7PIer954Wn8FMHAiwSSNI/qwuiHtIrASCL+Zfvsf2YrHjh4EulrCF
TL2owdibKR6V9u2sDp3YyimU21CZoNSx/+6Yf52/R2JfIRn493AXm57sz9Dk8MGyC6s1CBRLjgs1
2xmA3Kv08nMMx89C5G4rspUzxEeNzKeFukN1fo8kCCxI5CQ/r66rNEuWjHHLr4r72DX04NYeBdWR
PQmDqgV245yVpIZBP9gp7ipf7wBEMYZrYcg8G1Y0Wlu/pyfILa1FqfVyfJdkeiveMyRdPASHxUFT
K016yHjhArFV2xFkC/QiwxpFi9EvDrdJxVq5jgYtfBqxQNCL2dRXH44PSV2qKNuCaCd8KktJJwo/
k0dFnsHWIu0yEMCdh+ciFmK8RQyKgqP9FOxAEKOoUOl8rHuSEfbZDHhAcXqvH+WCxpJ/9+sgLixU
3cP0kTIJkVDQvCTcc4CdSZsj1r5Eog9mstrAOWZLMxzfgSSZMaqXlSlAVFWDcow7Xdp6tBbHKJFf
De0LP5KJYso8dAIrjeIpsNIWR9oIoR1sJdyvYzD6vnBNa0wHu6XCULr+/MM4nSygWCEyIkAV9iOt
Mmoyu3tuVL8QavxoJHJ04OAOQkr5tzBH7AFMqOB6gqOb6STbfB6WkEg43e2ew561EtHvfHMMJxqe
x1ziD7HeJUU6lZJGRboOmUwAJiQQPziuWMqauRczGj/GHVf1m47AjjBoAQMZNq814SOK26qPHhdg
gVa1XGuP73zx/t9LkVsxE9Mslvbh03E8wgsH5W708x/cXuPHcA4MDTVBGccacEsX0z4XE8CN7kyg
PcCkPBJhScOR4KNQwdVcEj5S9YiuWpQSnoDDc6uhH8AeDjWP5beDxZTmVRiHsGH4tspGttumjv9J
n38Rd2I4mDK3muMBkgZRGZ4OUZoixcNml2tgyA6kQ6GnBnO9bE1MLryLTI8Z4npFZUSCyIKSzfSx
hWx0g5b04dzfHtUFAlPGber1g/Ec7fsGuOSEDnc7M5Vuls0NcwltDfsNs8+KTalYe+lgs/3u6ezb
SGjZk6RPwpxSC23+9sEEOYLCOFucaTWy+0RiXjxqfPVB5Cl8dI4oiVB3udAG2HAFtnFr5saDVkSG
8OnloWflJBA6T5WRaUngs64nsSJQZ5SkFB2GSf0FYlC6bdmtNhZWNypoDcCnJ4jcdH8loLUHOBrP
V14Be52qa9YmugNGRLuBMZGyAtJ/95fDgqNkNpY93AVW9wmJgC+xkyS7Kp8ziCYW3s2jEHBqXN9N
VGdKnGmcUQdb0oIxQNHIoJW3UMDsqp2JVxcVdfINYb3UiJxj0cmcBOlIgqbqszyKl5iRQhPp32vt
O1wCAkGeoRp+CANcbIk6dLiYAPjsyg+tGeTHs4scJa3/OUnhE2vtH8LjrzWBRM2Z0nSQXtpzYCba
sQm8gsllssRtvAj21kWQCzGFU0cM7sB1ptVd9a/c1vDL+pd8YAxXJLWxBgUgnS3RakcU9J7p1CvE
HNKzKS23T4MFTJFjerV4zyWcf5BIeD2Mp7eyaDVIFsSyf3LBtpyR602UWyARjULaGWPG9c/VcXK9
xS0OTPAlqF7BNLnDpn6tOVmdLDesVaQ2BPK7r40z6sNQaH22ACMTFSi+cw9m3eeK1M9jk3Ffo4+8
M9CrJiDJBJffBcl+qKgZv+G5VZgBnyjZhz5oQL71vrvDmLdrJIcE/jKsnMwwgk9nBX/ATGEO7BF+
Vn7bMyk6vzXBIYseXQ+0Yr0G2tZNSSG7qR1hQYb2PywabScv/Ri9mB/49RNuK90nFyUuU82cwxDH
fQ+6UxCwweXpUCVi7uIbqJ8W3m1abp5A01FCoMHOZm3qXt3x5XMN04x0NkI67CKGmhBQwnOWhbLU
B9wFVT9ibKncGq0UlccCenzN3gr8CkU+rCIdyw9eM2iuD9VkVjDeetMUGo1UNVlxtVtHuglrZv+E
KaNvjmkEz8FKoC6ab/gCOX8g7NM7Az/RqkJg8Jz1Eeebm/RJWHCzqBnMg4mN/+q/OMPcr6LPXqvH
3tUSX/f5j/S7fcNBzQBDOo4gdIcSahaNMD8Mi8nfO+CNSRbYaT34SL9m+E4Uatw1sSXSUAQUfjoy
SUanBu7CGYFqElZqQUF7SyPOmfmAd8lJXsJYzyiJESCt9Qfp+UxtB/q15i1FiFl4ZRnA2zl87rCQ
NJTXsVLwKv+jSQPJsbnnI9r2mNgp7CCtolad3QXWbqDV67sKbz5/DOJgS2bTHYFkfpTwZMNXUF+0
TGSWXnMQg/IPjYi9kXgxKykVBrxxAhdXu5/vrXCLujfP2f0/R/L/w/iEc0lxgdpn6N7ahkFdunbf
bRoESls6baI37l44wlkrdnG6SUrDikNykH//HZ59pISfuqiFYw7fMwTS8D35FACrcAIaYhlVt7Cy
R0sd/hWt4fDJ+VxwA+bjt6T0HpSrYtkE2yNj6jeoBw7vOB50EGRrHJfMfVm3vbe4GeRuB4kO9tgM
MIQ0TLpMCXS/XJWqScg5ekQJUtbXNivSqiR1o0Hb2TM0zHWik61CgCyUGhbMgQxuXLLxHnrTcozl
lq97s7+npuWxzTvIzq47zsoma7GT0HctVCZp3f0f+9HHed/TGMatU0Zon7HZRiaoJmYwZoAdxY6W
dIN7kN7hvgFIs6prmzBeJdyCyfu2fH0iw1gdP4K0+QBNlcv/euEukxzSTYqeAZ2N6nuc+9/vtiTO
+MSDe9sbRKimNmFJZpzKe8T0i3w+8jOg/5KU97J6CTSW2RUoVy5w4Mbm8MhVPl2RrqViO7yb0r49
dF55oYxTMiVE2zsxz/9aTPzQzwuA+iqfIhGxaAuxxBqwrTKEIc32Y7f9mGm4i8/YcG/3Cffn1gwm
1s6kk7BsatXemnyulzUPEKhiWPOIYziF9Q8RPb54Z9gwX9nJv1DUWW8ovzGC/b+F9Dngqsy/9r2d
eFy3C59TQm0ebknkB+VClRt8NymfnNj7LnHF+Dnul62xdohtrFcmnX/WOX1eYUaVM+aCz1IqlaHD
Vm2EZtBsIOnwnYj2kF0vnrsclft99OPxrywWlE3lEmpGcGa+HLF6L23nzyQ6FJMlgXZyWCvcrs8L
kDjzd3mKawEWWQ1HuO1tXkn+pDybF17LTnTmS+zN/U/MhfgJxJScis4eT/UPS9mocIqPJfMKgnHJ
81Ta8iyGD9Q9Vh6T38LT3WFAV/TvLTs6zRrKRjBbP0ipPF2dg22mvS9CzEa+Cr5/VpqcdXDseICq
+0cHYp9F/5ZBUQcQtSLP/lN/lugE2KlzKph7Mx6TS5W8UQ1bxCrdXSxXDYb5j1V2UMcKnhfNBD6I
ZMRB1P5kMk3X1ffdmolnPQAPoGXeT+k5jueCgDFyCS+jI46IUyZEzt6noztq0PBJabyTh4Qrqayy
PcU2cXFdDu5FaSYFBxt797l50bEjcExKp79USxTsq0Pnum5jet+DnMQ+MR34yZ6CCPdW2rLlUqgg
JeC6ID80HEMFyApqTvR01HTf9XGQ9VUB+pmEOs3bftYx0glEdcqlqrfFmcWpOwpyXqkAwiRdo5Kd
nTR2DObh8II7r3sINo6PsTmVsNAUO//cmQU5XLwhl+K850v6nk9xWZYI14ownG+95YEYaSNZBYSD
uMtoqWj1EEjQ8U/8lod/Hm1f9PbAMYaWvc2equ6EF5KyDYgdAMLDbHWyrMOUoKio9xTSyq7YGDll
tzEf3/hwDIekKmwRECfOVpXm6MTZsbp/bTv5tmAtbbP35d6PZ7A/n5WHJmyZ7mcvLxfgJVKRGbO+
wQtA+rqsocovCNpqlIKiJvBXuB0Fb0XCeQQdDYM7kUh3Wi4u0GOsxMCvTfOioO8Nt04I/JxvtSsz
7TS+6LhVG+OkuLHzEuZYhNS31BQUHAvawq5BDkTJ7qbtoSIgyqyECNX0p3wlxlR/1uup2IdhVNED
shCBruWclLNl4OHm7yNDZ+CeDnfEhvDAc+ZDFM5lWeD5OpwTkU1uYm3xehwqPLuIfEuCUeigB1LK
6UDqtxGy6VM3YwRLTtc3yHoBmYCZMuOE6dYVtAfV8H5abd8g+9Ywp9dxLsZDF5QPxRv0dKHFZT7c
VIrAhIRFXJnypT9bnRqofzV650fRCno4dOn97d/OipXGacBFipTyfvw277/y1uPtObuYdkSorb8Z
zl+kET4Lp49Qmxu+RkU3XUbLIPj3RX7l8kb9y7ABA6O4S26mR1C+9sGt1HNwUBcN8p4KaG7UJxQT
cKr09gc0eoTGDraFc0v/dPdmbjObAjIHe6mztz2FCd9XL6CFPse6b62aVHfpRccwEswgjOFjeYKp
i+JAqeYlBIL4XE2wN7W0vUpUAOhOfUBoWYbpVZtS5kyG+52EIfYPsitv9JBC11u9YPgNZAfFIqAn
dsZNJlXqJZgZqvR00WJRTDHFjUe1Fpy70Ix0C/2+giHZz6QXZ2qi1awQxzozSV3L6wQdkPK1kUOf
10SUSzKB9PhsxN7r0aw94zXpqNkDGAGdNUGU7ZKhj8FIUjoUmo0c84GOx6JMh6s9KICrqssuDhHX
/2GUS8CztmshIeQv+kqtHiO2H6Dbv7NNVUWbprhXT6eTAKxwMd//nOjuyzvJmeXPOHh69ma2LvFd
cLXoiY038fXzflG3DHTyiqDVRXrsA+DjCfIB+4ee0V9JGqdF7SvSZ0YIwpiLvhia0Igu4BHvD39/
+YbFWIjX6kGlDwBPeQFNCrVK3KuZoezUHbBq6MZsHQT7kgdFPPhT8uHFTFY0xLMeNgODs9s3Wq0H
rMrUPKaSUbjh4OgfjLbYg51xpeQLCT1zcAEEByM8NRQhfgdpfqHdd2Cf+i39TyG7jg8hrJ7TFPiL
oMPa8EmxCXnZqa4M5GWHvYLa91u7w2J6/Cg6CjR/E8Q/E/uiKqMkUuQD3UZjq2QWlUdW0IflU32F
4T3U3BbACso5ts3UvT5m91ajahmEn+OgL7T8TM+ntG6RKhSargEblENTzZWorBqNJ8J7gFJCMp4e
ZYnFjyDgsIaXBk5f4DVsNvIh6MoVqy0jnztC6M5fB2stk8JSGrWoPbzoGmqaRIx2iw9lam1GDajY
AVcjAg5TbDraKHjXmJRUnB1BngOQFPm4BeXDQQfq6kEsMOxrgfjvf/jdDoGrsIZzG5D39Qgq1LqJ
rrgN530b2wxh0w+FbP2HzgsONrO1fSF4TCAull1mN1DHoWhTWNpcathqLZ7ajWNU70r6nJny/dBk
7sdn3a62HDLUIq2kwVnN0ziufeKhszv/T24/6hyICTeqCRKIb9pf1zQs2f7h1MIQpkm8hgojHpTt
cz5eAL3JZOMhCgAGgsIuUsrvOgMAbEUiuMhUJy4Nnpbfd7m9rRLn1BWULjWP9Bdy0eYyo2jxX5AW
tMuWoBEy/hzCh9CPHwAJcxAOaJB5sXm69Ny8fF11qOwVIfoj5J3mHhkvk4UOAArBY4+hfFoNQqIm
rrrO2mhDc/DzHwxiw6HpBJIkRZSLRnZN6rsL/qjtaVPKqQhWvGEfLEc9Uuopm+KLn6yhpwyOmE7C
7T5ZORIm587O8bwJNQX3bzE1g+To1eUQsnnX5LkAyayM6qxhQ6eqMeXlkpNoJEl+I1WiaC6TMb2O
2LEc9DJ9mn874gk9kRuRkBGtdox+yPLSYjRf2+dPtKa1lw3e5I5l4P/FKjQ4AbL6P85JuHubJwK7
FV6IUdUo4eMQtHR0Bb7H1VBuEC7C9Pbwu2UTi0zI5cTtlYEoztctzA+6XWx8qMwyomLqfjnmUn8N
+qBSBcwyGOBMln/iX3uXWXxqrtO+r0y8fXOuMExLnyGdPY8unGkCnXlJINhPCxHvJd5wc55CNpWZ
CBtq0T1tugKprfsVDVWq3NEiVDzjJQyyEhsyXb2tjCOdcB6+SCWDXY1Jevs2lavz/nfza0/iZO/N
gvRZcnHlrt4RphHENRpmh6mLTRaJgaD14DhsElL0VRfaj/24GdIeRalCm72WD9LT5BSJHET5645k
tvjLG8rlcnXNirq3nJNMShOEyJy5rl4wCS2g34ypkADzyNwEeGXA1TAybYrzQ3FwvznLNeEHyWy1
sfqwu6gG0GQWSZaZNKC1RB5Rgi5zSua4FyD0XhDIO3VHSTrtBZs8ywuY5Bzzzsj8Pt/CQ4wHXkNi
5YxWMrmHWNcepNKCsPa12ljzm/qfTgATCGl0pXrfzFFuftJz1alFFvqSZdae3fTdiL3TelxukVPV
qDL3jvrSKTdYD8+T+XYZovCkoerhcioCHNB9v08qxCAP/kd4maotYBQbiwvn1pE1ucEoGflwsxOH
FYs/ckX9XHAB45Ly36+CA98vid7C5LbtY3IJTVYIyc9U3Vrn/EIvb7ZlaGBz65m3pK1FmY6xy0yo
1ZW/cvXHS1if6c8XpdtQ8Kpi+aZHpZDxqpttSsuzaWCF3myYEKlRunkEwQYVECK9xFodhKTk12o+
2JGDgLHcQb6sZMsCSx6WfojjUdzzYyde9c4kRUFK83AICDpjbRMXI8ZT8L0bwI8e6e3EIWgXBd3I
0xbhrIgXda7Rsyf7NFPPxu18bwNw1yntC1SaQe54eVRlASQvDLs4duQmWEfUjzR+WQpE6ymV0lP8
VAVuFny90MI252YmraFYdhGkw3hzBF/uNBuyomyMlWFNdvbTGhkiJr4KAazyuuysro2CMCz5R/bk
JXRCuYK553TOjmIU2zkXu031bjs0bcZn9mbfr3+us0GJu572Tp26zPlqUQgFQd1OH5dp9S+0kZVW
2sF4vtsIVNMvfNHRQMBtZvRURsIb3gafsgaySGFYYqeg8jUSyZn8xQ9GK7EpBuF5u+K5JNX4d5A9
xMeeRhdj1TR/3/gxw5lbdzFzuavA9cBJlMWzt0v1iD4cYsIjj+IecPitSM5NG8EAlw1qcMQ5/5bE
H85AFb5Qnpva0sbcOuLnmTqOsyHP2gv0pjy0zEeQ408YmsqgH9RpfmsnHUXqchu7GhFc8vaw39ET
Y7ufLK3GOz9pkvf/76mCyqm1kzjbBwrwvc2MnFevWRUaKxmJSo5Edyp0v/CMOX+Bz/MbHuI0N9AX
EZdGiSIEYJTuZzGp7xtM/BZhM/yo1s1lOuadiY+lzx081vUQ0Ja/zKcY+2DNkEoWdMrAaX+Tm2qy
y7wGHM+X0tPwCXzvSFuQLvYciqx/utVK5KGLpaekremAUUDDcSbwTYk4j1IMGdr73/hqgvsQ1kBP
B/mBMfbwSbE6Gl5T2XMBeFuWVH+bEzDldBYn4fCtuktO2mr3LlZG89uK+pRCgaDKx1nZE+TGURRW
xbO2wu9cArIzzZdMWj5/xKRa5CgsV7qXanUGRa6R0E+8vCFhJ9oO5pyKOOkPsxiQDxo/+Q1YwUay
LUQcp9CLgJLtt5RfUiA0cO2SsZarhjxZObEUBp50JJFCu4qRgDMCb8eKeLrsA2/h+HUh0io8xZc3
8Jq/k55C60FYzZMBjTKHjYSOJEoF1YV+yzHz/wPfXq6MS+rQWQs/InuNvbKhm3QTDQbruATl68WP
+wxn8vT/xQS0yTLW95rufpbIj8FlyMOHp+dvkKfRlWfsZhDNZEoNahgnbDbQ9fQEw0y7hQPr5+PM
kCnGdC50dDD0sic+3EUH/ELo0yNQ+Is9aKSu7kRD7zvrb4KFHG+RFNHoN8JraeGy+clB4TwKQZrV
kiiYrPFtxwwnIAAJuAEwG8GUiGI0gmbaoJ3yeqIVKcButsEkEvLTGW9K6HYm4/mdcdMIlrmY4v2/
uSDUhm5qdWjIWhlnE+U7ZZVBqZysa+dS0EC5giLgVtEloE7/Jx3r2OccpU7WZOYAu7T1lKlYrvyq
FuO/hRpH/grwzTwJqHW18ciSasG21ZDHIULXfLvel6MIn1k2APahIl4qtmdGX5V9ioDRVcLn3ySi
YylSeUujI24Hz/KsRTKHzreMOkHTx5CDL3eVPXIthKObDxC3CedIReIZrSkXH6bxg/XNTISy8/rI
+KiOkuDSwVT+5QOMBNRho7+fx1AXmnfQ9N0IdUibzhagB1RqSE2e0y4y4eYKlz6p4Fhrw2HqkTTX
5m9zjIIVSrDWjEPmHHBustPB6v82awC3FXTNDrkRGpNgpQsRLC0BenECGAuXJjfpWERPzwIa0zSW
jNjfaNqP9BeoVrnmH1zg0DIonVnWjV7k6KtFKczyhfigTfN8KUOJgUbXdchB2HgUYwSnpiXI2KXR
KW0dKKPJ0DptiSNsECHMbpoh283GmUfnW2vkx1aVLRr7qG2q8b/DO4u9/yQ41bk4bK9pW9Ckmlde
V2t0kwLVn5tnbhvsp53xsa6GOQjftIPHqdXis/+Xi8zULR+ZyctAj9xaQSOt7Ut2Ba5zbReqc2xq
K2gTJC0f9Vft1btrTKz4YhDzJhgb+6xFiHy5ENuthehNUZJj+MdYCPKBB52zceAL93Y8nwfaPg3H
XQtJIgTIsZdEV1HVJCzmmNfzOh1Psz+soUwJpe505Ku77XzSV22pam69cKwnOacqqrDWA7AucKxV
IBOenqV5gtchyKcOEHnNz+Q8I5mrW6iLk67blYwy0UPegVUDshspc/5rLsXUcxuby9pIeH9BV2LX
7Rr6WrF7sypi2jvOY7YP8U53xzJTQ9xHcNC/0orBfMNy9Y0m31nLXRK2eBNRE52Mfrz+PXTOfhx4
TbCr/op82FbXjXL4PwDLvweVMovuY/dWQKo1ASFAdxmBl/QNiOYVtdcG7mDdI1lZOgI2TyemuuXn
2Ell7PLXuSSUuTdvaw6mh62XvPZFgOMVNq4KjjRp+i0o4dek4plt77mn9hn7O/Ods+p/Pwbvy3qb
8QYmTVCLnBN5dMSV/OtNcmOHhBXioJiuUGjzh02Jv+1OiN7E7bjGdyRPlevxBL+Q4xF0bL3zL393
zQUGBv6dHGIRvKhYWsDvI7B/o/fCMcnwStvC6mP9FzOD4aEW51ZXaM/geKhK6b3zDA6PYadLktu8
1G1QO8/93FJ/qiujm/MPJDVfR3W/PXn1cFdu0zvlboTEVYD/jFWvradrTkbglX3C2PN76UHI+JS/
jQ91Lhqc6xxpIO325IADb696CsyfW20r4JFSJSGLhEJlcsoUYXGEogeV5liGyrerZbfhhZipH+WV
9XnpaepSzXPW8aM4usl3eEqEqNkyWUCquf0+usE50AD+F8bc+74dRzhREPCpF2qCghIf/6KLVvDl
Q+sKJDt0wAatdR5gJoszLfl+hmhA/dEeBmc61tuwAQ7VbjWQzU6l+iWam04OO/sjbUC7pDRt4AAe
q1D3QAqRTrMncq9VPTykghb2JH6lBjNh9asx9Nd5J9pPaMYi8QjcTPctmduDRojAxZP+k8VZ3UmR
OBO+D/ghJWIWiTGiZ+6svWVVIBL7phNHDE65VQz1SftArxweR4XxDZJapJGhqh8bvdCp0z+dx+P3
nCxbNQhNIMD6Zah8Snht5sEbAFOeWD3l8dJaFYHRu1aQGMW6raTxdR2S5ubsCq8gGXr7S2Kck7ZL
TNbUNU9tlWwWlMsBWktPPp+wHVySMKxF9ISbXRSKXl9uUVIerA1N8EYSA1yYcrua1Yvj2+kPqAQh
13EV3YgypR96JEbnocF9lELXoiN4hN1LPO9673lCTtwhlEhjjghkjOYjDo+0Lx08kUu5P8HEcFiL
Kz2DUV5qgZmwuWtwpEmfAuWsUTfXhSLx+SEuOTYe/UsnTt3XUinWfLLeEbqeVPPGrM/EW6W2Qagr
SAcAe1LX5XY0mBDHEDAGy+TcKFDrHxXEfw6zjHoraNoJp7aIS8hCkncVsfPIZy0C/asuBzuJWgRn
juVVIn6WBtyI8Oe3TDElGPnWDeuzRDO4YXR327a62KeobeVPba0EOYNuzcvbjiw8nFPEkiYtXQTB
QVeqd+1X/GNdyImU7TFOCqOW9tpSUsVuh3wUrE9B8Ad5e4RYe7VQZTCtWYyX1HjzrlkLI2CwDJYV
r46lcGb7DdcE1AcBZi4pjLo5VxFDK9rCkEebtOsUwqfkz2qR6vzO02pjgcZNIzWBfxWaaDhKvON+
LOl48xBO7ouRN/YHrEY3LwkTA1W4V5YVY8GoLcZMN/YphhIdkX9MjOgPXoBArycJqWr+iv4ECnjq
jKsxE6KzM0WdryBrJrPOBKVOT/JPLQ0zsgDteD7ap0THyp+c7meWxAch2GShJ8qgi3HqSQH7W6DR
I9p/+tlmbWdapJavZoId4Y62NG+/TRBEv2O1qR9G8fXUD3YpilA5sfkXrJI2sF/pXQSX2bZLRiGG
HFvs4dGrCbfGiSc4LYjNqz31zEwg61ITzLt4kKd0DzRQcYofzv41MqtAAVpj6UWBZTevjO+ZiB2G
U3RYcH1tmoLihu2Zg3L2NS/whmN94abGnNWomEy+epUmFS3TJwZE+K1UmcCZSxuwIhDRwVpt41R9
m8t7QQvHSGOOAlqCqm6NhORje9CFtAgAkdIdTzwypQ1HMBen+6wWdrZyTw8fmVN3t5DH3qaBH9dL
edMdV6XZiNhmbf+E46KxBxiarSf9Wm8VKedaSG/EzgF4XAXsvSMUvVtLHkjCCxD5jwtAEuENB3DY
VMY9k/nAg3zdDTtq/Cv3VWsDb8jGD0NZJmj4v7R8kzqXn0BIeSDKr539bFbtVTfv0qeWi6rasUHS
kF0s//Z7Adh6tTwe3RqJBbmiCjzrA7zqyiqjIV1Ld4y+visWTLSvHXEP1LqFQPbC/sSXlO2jdaMZ
/wxeZng/Eo5v9sehVvMLEoQVzCEzxWxORoBjo2ygTfE9YUZjDshcVgVV+FaB1iwJPDjfZVOHE2kB
dQhONul893HevbEzgIA249RrvAsmCq9wTItlPwqEiPZVrOqWcXAieafRYcj4FlYBIazZe0ZA7hfP
/OlN10eoCWrlctoZgjMIytJOLwrifoH/1l54RNR9g7JZDCcPxpbaLwH7D1sFNjwsbLl/VwSm5NAr
szdOSQzP3DiTXPV4G84q0ZFS09tIzWOYhWb9d8ATxVrNPKg+yGXJ9WLbq/uZ0hpuJGaW2RU7XgOJ
vfR3hY5m5+eCUJOgsND/GNTpqEMLzzuqxrf8SqLf5ZqmVd2TapiDizuBtyyKwKNbiB7RBJ6HNAj4
f8uOzIQhrCDKZwdshV4k8A6KF4S6DUh7Jkigq9qrxFO3+UCWtkjrsirAA3F4uwWmRZuaoMbhxbJl
+Br4DXMIV7/6nLDDrUt4g7m/go0tR/Z3KwaWv14VsviyaAyCfF/+CVHh4gUn5HUc7actfR6j3Mgc
gp7DpFxE5qJd4eK2VtVUTvXDRGBH/vpQK3wvgW9BseOHYAK38uusuCuJmcE77JBMZt54IMhvSCTv
XeXLoITv5hmcADWpw+CP2YHru6gPFAXtQHXiPIjhtkH2Cdpv4vjpCKzw86r67HRX6nJKp8pitP+p
R9IaTA4wi7tUBNtctJihOpTjrk6CmmhVs2b607k9LxMBXX74kESlg6QUSsjVX5YePhvW9eWhbpSY
CMemSX2eGc8Sfu2jk6yDyaCYWRuSkw7zWAHMjIIIZYz3xVdy3WmE9vcGvae8tNtxf6EL3JOQoQH5
oip588r6LAGDKxepYcHW3vfqZWZFn/VqsmR6cmxlvzudHBzrlHh0XJ8ANKtTKPGN/rp5/VE5QA8Y
iJC7gS2UGUmXYRb6TEUTvzT7egdSTXlPugeP0nb/7RoiNgG0ffqUgTVNh34+/5WbWoYPSoTpz26m
h6WfBAQeq/o91SU9wMbKD1YJkM4WklmvbHvj1NU22TDdh3Blg5NqjHgl6l2HbHdEdLapB4Nr/ejS
6ydOdDn/qmk3OllkMmC/YmaoqT9C/Y4w2plKD5ew20FLlIvRPQYpH+rmmfoBLk/myWMVLSRz0MV/
YwbmXU/L2VIYCld9/v/KwpH5CJTTR2XioswddrsZCDR89UWHadAYLwBKadiCj0y47yR/RR1myqDx
ivBbcL1JLgrj/fg6V5fDXQ0UgTkhNT5pLg1NhPiaCmf4rVL/NCIuloYtfMVDBvq+AjfreIVOTEU8
na2hhTipJHBgrIVjU6EEqqsQC1fURnkzIBQKVwxG8lqqSP4P9SEKeL1n9kbccX8FGoIqwK3WhZHn
/iB4G4KjkSfIAIoDrZKScDWTrOfC5s3DJiHb/2ATawO52w0rBNUbg6yKh8of+Gv6MGLtD3f5Bd/j
8axmplmqn9hD0GmfdOtG7Whh7MAfNVs0JcGT7B1G8xnNMQiJU/LCcG57vLd8Fi4VODXvXJhUMyo+
TsC4F/DA14bTGpA2K88Luir/L+EJHK+zF25913KqXbbJ6zv/vGvyxZZfUEJnoS0I6VnR76qmu2fC
BFJZk1ZSINVWytaOOmr7gLjNt+Irxkp3oWpdcnvALnKOU5P4C4Cn+pl+9NQ/flaHblPC6z0nxw6V
zc9CB/GPkZqqpXnC6iQ51XjOoChhmZlcIcV1vMtgR4I6SHhcXbbHXC+h6pZHN5JRl+2cCRMQM3TZ
owG0LMDABTEG03gUATiIhj5SMNL+EevhlUKI5Xz58xLmfX+M9/jbSBmxXwIPuCXO3EKsE/bB7xd9
yRjLjotUtRY4sioTbrgMxIpoFl8naATU2B+povwL72bXxrxJ6ni3+vhtxEg5z4nwrU/d0MlWmD3V
InmPQRYBZTwFj80ARj2KasLz6DhR9WnBRZqRvpzHxWEv7/R865qbouq0oayn+BG87FLlZkdo4RCR
cjyFVRQMVlLjxsPxe/iMZYtTCkayTQq0hF7hHdvvFAq/ZI0KOJSihK/7dHeIIy2/EZkTgakJTCI5
zFRwyq1QYlK/qMlKLXuHZm+EhNhJ/LsP1K6GDp0+M+/zgw7ACQjaJikRLKn1Xxz885ozCvjPkpQd
DPpAeoksfpSMSBjRw4iYXOdM0t2PhHTDnYXeceTGpxtCv8alHb/ddkXrfW96ncqSWbgSLhAcAX3/
7ghsWZ8HFa6sxu5GlFjYKeIcsZiRmqLG3bBC33TOoXvL6lmpJC/1te1QgEsKGABRNRkKyieAAxCV
ucHA8wjRTUkqg7m+fLriIwFWvUq3DW+dg7Kb1xRBKl+zXW9iJ7/jD+WDBUvtZZpfxAt3SVkmSRh0
PbDY+Gop8rHHq4PqPPJSPDDcoXvAPYe1PnCV6y+lvSi5ZWEqi4Ev10aAUhqbt/t8oxPT9RXduq+D
xquXKeveTYGbk7lpNcQYLJL1gy6Re5jrTEQjbdkbgmskoYeei0guwyQUUykxfhA9/PnRzL2C5RNz
yaCHYulwLSEB/gz4NgxeEDzEaElD3u/Rq6FdfqdClONeigVWreuC7p6LZVZ3JGcwUT21xx/Um3hu
i6+CLQG6R0QvMQC0P8nnFQpz5GdOff+zrkZ9PQPjw1f35iqEcp3Kfxxx3draIx4KJ+7qUzaBLegN
zzZ+TRvv2gIHUbSw2pL41AmBfGk2R1QNllIyCCR4thK4Rb/lXnvJ3+UBpjx1i3/MIWTucORsUkVQ
VbPehWPAjjoL6JQBZj1I5zOoeTzZLzDW+sGK2xOiBUYO6yDICSLeNnsyQ8xoTt5eyoOEyJLSXyTu
CUTrVRypJe3/u0mI9ME8PZn9zsAXfAHcr/X2kSZUbQ5hedZF8QZfmOCP6+CAEWun9oEv63AfFZ1X
bptLTYxHVaaIqORFrdgNtC7axoWTpXHhyje3cAIFA5tVEogwWXPH117iZSMHE9afmFmZAauP83k1
VMABti6BRdLyosDGvI9lE+0LQx5qPfJTEBSn+S3LA3z2z0oZnuMBFQOZBA9vkJSi89p1iWLhUC/E
xzw5lESwCo3f/X3/42cHll3rbMUOkYvbr68SlbB0KJbOhNvlRW4kliGWqRhmhlgO4X7842tt9hM7
qoGxihdyp1cfhgPIjeIu0PmT9jxwjS3afK+P6WGKyvSnxvBnriPzX2uhaBfP79Rfw5wrFLHx8mr7
yMP57tl5VtpUS7hK5Nkn4rpHhJfhV8wnKi1PMiM984URQGGX5GquL5PtiFDKjzKJ33GcgwtpE2aI
uP20nh0JM2i53YO3Or3NCctWAAC8YpMj2/cy15hTH71cyCOb1e6l2dtEBhhKLP+X+AGiGnUJDlQq
IZ1EGGoc3ElpwG34sTGHfJDk6nvP8nPvm1hNJM8LCXXW1dDznxHLVYCjHTcVJpymXGeVzoVDHsI1
FHwwPpn6LIZCkfVYSM+59JquYyFgTLlKkXPx/GcfSDdIcIZkFZH+q6sN/2wPq+nYoV0p7orE2GpB
hABjsHusJh5lF8O9W9uYhzNDw2CE16RzugzFGq08F+POXr2vUY3J/yBOgnneqRJcd+lFVbmoQljO
kacePCCT6s0gpeSQhNqIOKfpqxbEruPT4WWcO5XffJQBVvmzRFGs1AsLQA/9Yl4VAf5TmEbwFqgs
K/fX+iuKXdk2dww98B1BtlK+hFSQIcuCQQP3iUaCDmJrG8DPiEwYzUZJxieJQxCJ9g7G8GVOOQrS
V8/F6SCHqX3VFxCDE8TWPj8VctNSXevIqbz1M8iiJXxv1lr7nsmY0gqwMbrgd6SSfumjCaiQElFt
sLWFsAOL0rBhdqyIZ+woJULu031Icm1l+FMVz/hq3iKLWV3m3oAP5bRjWjWPI1RfBFKVa1nSSw9W
bQs+bUTNUBr83htMBhw38/fIvZGXpuVZPukzOBH5bLEvpAvp+1Lsoot0GyAWq30Jb8ClvXnCjX11
+UhSBgi0M36sT3+CIenZ/fgtgO3aHH86BNI/w79PQoAPh2H9Yp2i56+X1Om/UdaeuslWKcM+3Oji
mpihSplnPsjHQxsExezxmSA6+I/VImFFxG064FBIZcptjz9eFqw8JwK9fWx6xC6Bd1lkzTvNqHZl
oHT/Em8BYWxU+dznnYr8h+a8+KIl2V6bHQU+oEbtkvtYOeuSu7BgNmc57MicuEYhlrL1dRHcTaRJ
a2u3B6sdaeJ7YKQg4XMzhMweMThVvMX3BwaQ4oG26QAemwgGNZiHKBX8zan8BNBKQzqi5CNMP/5I
TqOvI2IIuIRRQCDvsA1XnwDrtV7eos7jLHkltUxW581Fl75avM5qEiAAjMxrIrFxfYuRco/ZzbDi
sdiNfJh3yDkTHqgfKZ3pj7tAi1Y+D4lcRruMXPrFWTt0z5z4RyRmcQIyQN0mlqoSk1XPJ1YR64Zh
9hXC6C5IDwIPPyNsryiySHEHEZeKvV7P2jA6upuB9uw01CfKh6j28GmzaHNpfDTvM6wdyMj2oLqR
vrhvftY1JOv/X393eEGwltz1EQSGHJny/5+nMQnlBOE6HYcDsLTaYhOeybTvaZTvMrLFi8w5Yc6N
3RwntDeGDnCVcnRQ1r4mBn/lzl69F7YBtwYd0zjAW2mITllSxmZktCkaPoopxg8OF7ZHsx84JSDO
aH5yWKRx1wtMBLH6nv3vdpW57vo2027NNFu+j2TpHUV6AVqCQZoD4BTWaDj2ihpEL02Skx/viI3A
BR85WHNcATU48ZsW/E5QsQmPGlAgVmFp8ybeBup5mBJYzpjqj6kWXqAAtPsTcAjlbX7aNR4sisWK
6LTCDZ9FdRdZ9AC8VUJNGRmKvvhVojSSxoRrSazrQgPeQI0OQvqZRoFZZTHjQASydLdjch1YyZ7b
98NXejuv/L/JS3qnrEQPPvKNys9YGgfme7R1g0hXMY1XnbAVDEFkjR+NIQTLIxSLgIhj+gI2RZ/C
1J6egAFfC4hKuOLirs7fwpQ9S9DQH5tzzirNPBzQal8IsAzKPClbNTTG+O0+SbS+DAy99IaToiUj
osyta/qwskm4R+H1+Vz4QPqJnlEJUOGfOuL9v2DL9+UCIBAfCCxz42kz3RN3Hqzbr3pC7TeEVDZ7
6KEnkHq90BPu1DNgLCitYmGNkvFs410uZOelAEA83FYwshn0iwTxUSuWkgq0IHcTfv0DPhZP3641
AVRf0pNDKwkE6ehkBOHoxbp9+QJYtagmqixCOWa2uMTcpu/rLlrYBcKggmBZvc0foFIKpLAhLu4c
kQhpYsaZx+v1aNjTYlvV2lilCKppb69Ken5U9P3bFwxJpE9ABZvqyeoLL+zsN86J8DRF6I6AN6iD
kXb/nOnlGj6MPP8esDyc+/70F4AogqI3uGJy8UuGsKQ6G0OMvJzoS3fuxA4D6YHTLl54CraC09J2
H5CaClAfDLg/rcDLL+1QGFeFjew9MPzzKbWs1sioBqUvQbwWc5ItyNz4+f3zH90Pwol5lhMyUflW
5A3rX1noLlm2jY6vPKsnzL8dwBcy08Aq0joM5HhoQeyJV+qMm5jy3uiiaY+vUm90Px3wHW7IUvFG
qMseOZW9PvoGGW/6aiwflsC4/LXOstcexG/g+6RF3lH4wCymzoV5tQZVoLH7hmd8mDf9dsXPFR3p
j6dRC3JR396VNKegf+hVVM9GWSqY/UGnXl8wbD0IOPyqiklG9olXUPy3lju5QQl2m924nLlIxgA2
iUSPepQbbxkdi+IUV8+Np9SRpCku8zzTeOCwZ8gfgtSWASJE4TSVfZLzjccBEMCynuMJR1rGcUXB
d9lcJJ93B3GPouUVLIY6rl+kTFyHGZsqeSmeg7YdaBVYVSlaEkr9gnWruk5WWrxz4O8ZF1TO7DzZ
cfzdzckzaxapDXwYVe4w7LJ6j2pUqoOpXvwrHzUALSwR6m2i7anaftipjFdiGjdK6ZjTYdqwEoAQ
JW7BDGX0QPe1B3mbZlAzJqZm3O+F9zFDgtTjWQCkoRbiWka4qFM0RG41uIs0P1Y8xa3M2eIH/Ytu
nNXfOrEtzoE4bJed8gxxbuLDw17DscJWE5f6r8rAWzW2Rb9ymSI5gOR5GRSscxyOM87s+Mo7E77l
3GvmeH9zionh2YGa1rxuzO3aaUKvwrXVO+TJ9fTUTV/HDdooyPpZJInA+Iu3mUh+mz5S+0no3BiO
9lnMEjyBl6Woxo8D/SZAJ9EEpVC+vDOBY7wuMra2fgvT9IMWVE2C2IKER0HaaqmPD/W3e6/f1MRj
yOO+3Toub5Z2kqT0TNNIDET7eRJ+fHmQffVLfrM+aRyLhIwJ3IiAGAlPOfHbM2ejrqp/3wIwjv0D
lAY4s8yakY5G8i/bxFNLkXhEI05Om7mSbbhNnjoPi7O7D7AmCT/wTyDhQWtMoQvQHkg3xwdGYwCW
zdn7PmTCkjxBFJB2HUy5dqIvSJV/MEeU7MnRcNY5/+wyQn/hJvo6VCf0gJTyCiu2CHWLBhKW0X4e
M3GcXoXeLxgq6HPJnsNg8+0Ga84YC05Ncz8Tbao1jpv+OtRZVI04V8ezZlqGd9x6A8UaIP93DFZu
tBO90Sqv/YYIynnBLgiyRNj13zmg2+qtbxEiQhzL7fH/k+8+05IHWL+SLo/bBBydCe03joDBXEdE
dxDpUE119SZGijQ7EGtpAAkdU9hq4X0PrWnIDWo/5S4RABJ35sUXXmzR/xvsT/EYlnT2OYgTQcF+
zP3gvbMVVAIynBGl4Xly5RrR9tO+MP8SCqqjlJizUL7Fb3aqsC75+RFR+/gAHHEW6Emtd+3poei9
Qm1fO9Mmyxp/vSMenfpDWD2ft+jbHeNQsNb0Fpn4Fm9CdRtW9TwzaxAY4jyi8p82xW2yIkvhWrLH
X6638Q/VFDxK9Pr1GB3PIN9e991QuinBc09mkRNBUJPFYGlO8nVFo/7X/084K4psANfRo0B5xgqW
zp+88uWMs96K0dx0V2aYUEL8+U2843XNF+BD70FuEQcYn7AYC/2fTaJJgbqRm1CiVvAYdS1zUiBw
b5OtZDHD3NYY7KbLAxvDYDhIETiNufNxHnuJiHX/peqltOskza4WJqJ7cL4yo8u2tiVJ+lFlwQb9
hiD9oo1DuNBUr8aOMdxCR6eMwiKqMdqiRW+DQHJdXSu5WnX3d9nxg4EFNBNurSxx83UustuzILPR
ifcK2uoD3QcMsDAnlShO/52eAvxVzdq8JvatInsI/IFzJ0aZr3K4liGedzAbTUFUXzgrutME/8In
aUqbTbKlapf+zFVo4b8t7zvZnf+mH/8Xgd2ApiBL1HirCUJVIQDdDo2w0nfaPiHvXqXZ3ab8Pgj5
TG/ulzcdTIaxUcR79MFeUNELiD2um8qpCSxErhtl6apHxNEEyeJ8rlABSYAemNxE6frN6txA1iPU
+CjxNvp9NrqUjLYgsF+pAAwoQO9UvN7slgIDUPcZ/EUr1LDWBE6341in9hhBErtdE61LIdj0O0zO
VRunn5ooZV92kwpFCCPTEbncoVfp4VAysXIG8gxdmvXmAwU9k0GgwBbUp/yBhMndmuCIeUszkFvl
lN1f458eT2czoro4vG/46vIfktzPyteUurbruU751dior2zYEFGWoNwGkeA9/nHNni+fNNbjIvSQ
nvdf+k0f84lPWpmnO26OgEKOLnCKNbgCW99zBxJ0F/Wf28bao4QEauJnAnPKki7g5srdQNAhvh5+
sEmjOJI4fm15YvxgHHHAfLoiWVSdw0tJ4w1//kFyaSsLkaImVOT6qkIj1Me417cMXkWzLi1qmIh6
eVR9Bv2OLXUIxqCYbWoNtW03D752qSHeg1sTvBcRkDI0JRSTYIhY2v5l/uyJSOCKpOs0PyrOZcbm
znSGIUVgX8aIwqIajlkQKNLD4EWS22xa3yHKIlG7zULdEsOMQNlBrezWZ16oNGkr1Kcvgis34N2N
d6O4dZ5SC8I6KgD2QItrm6TcEEOnQfpal50cCQtg0PE65d5WBEJ4AA1W0tLyTc5uZkECdKPdWLi/
YgIuro87BgxlfZP4D3Rf8wEgjxRkOcDuDOYRsLj3o25ysbVC0Al+9wDKZ3YXSc9cLFmFynrIjsd2
pOxfRoQz1rU/uyEQVqp2rgGqerRmtWyeF7PYMaB7PDLrorEOIes8vNijTeSLcqyXVutgOW9W/ynV
7rIPJHfBbxiSK95jGFLL4NGMe2L8X3KoUnWKxg+2JMKWC3drAjB9zYyTcqRwlgxImKiSlNMFBcg0
VW9e2xe9aQDWYpI5dZVtk9LSRYGRdtmHR05EvSN1YsZszKTovUfzUIgQlpH59AHXt1UPROZ/K67/
MyGyuWLR7JsJr/9ONGI4mjgFF0bn/O2lT9Qpdq8cD4QpDmml0fRH7sYznlMhJdBfGVcnYoR9QDNw
iVpYYvPkvjhM25ncACNZls8svwuGO9A6xmsQGbWZhh7P1F4rv5lujeMO/fp527QfOcfqGQMDb2qr
UmF1VuZPZKYB6A9U6dvDwPG3PeEbuQaYJBq9z8PxiY1uYkt4o/oUPIY9rcYB9ucZRIR+N3i2kCrE
OE6SqLVRwWCji4jfji2F9mqIWdgPxljoaQyCzQg+RXV0EcG8Z3PL0nRTPVIixtxTSBLNT4rnrLpL
p69CLM92QuMqlANavksGKSv7C3PKu2hS9dZc9NTC7Q5M0mkMQrKumZGkbaPHOpjGzRWMdRocmp4U
lfblyJ3+o9ihGOLKgIYs4nPoFclykNqEDsXyxq26MNcxfBmeVSZuW+SDE81k1QD26Qequc2LInZZ
Q2YwtVWhTjZyZ5lB+jlUMhprUAnF+61goEWx7LmWI16KL15uy4fR0yuSMb8s8LD4oRIVz5QOsEQP
2fSI7iyDTm8PSIYkvO703vUsRC+AbriDJReckQ9vZEnwRswSDrAYoAMHxT8ua/w+7KJwxfIZ93YU
+vyE6+oK9haxhYYrP01j9V9m7HAekGgU6yT6w1mUH3DKkJy/YRjtiW5I/strdZ5/D3BNqRoA5oBb
odswdZD2sjZd30jKOOoSd056Psr48pHR14SVwP8y4UKpjxVK8mhQ5PCeuWtAm39p8jSX4LpFAzot
vt4OgGOD7ePoFsAmbK+cnUZLJIFp3OFVcTpjdZyd3wivAUL6eMAJdsTlVmWDVQmz8bmobb7vXxN+
L9/YHvrmclstXo35wSbhmoCa+ohn46oNaRRsHNuGuJotcuYfYqUaRZ07TdDGiSu6ptwaKF/1pl2o
+NqRrMfzhog5WaJdqAYCmLrweYLCn93kS/qrgcY+wV2zk+AurofNUw0fdfEOK/Kc2Yi+1wYOtaZq
4dcXRHp5y+ge3ySOujdt+uuwoo+6mJKHf45Qn2a8ZY9bKlpVeCg4jdbWXoDkDJmAi8tTZHplza4x
mV8QSyxX1W2JFigh+63kWk8KPJ9Dd+ZQO43BJnn8qsW5zV+epTdBLqIRVxef/2lfiQZA2NNrB4s2
3TKqrA2bjbKD0dmO2yLONszgFBc1RUqadED65xVlUpQE/IPTCEf85AeOeMzD1IVnnhDg5beLJHJ1
7/z5CjzGGcO8IDa27rexSJKIrOTuuOOMJ0Zk8yDfh9Crj3bZ91ahtyhqCXWqtpDjIu0OyfNGae6R
1LUkyEpce2Hmv+RYgSlWZIUcIPkdiBYm8IGaO/sCaVS1xZOtHDl2Imi68DsIK/Un3QnsOi3kNmhi
5RHNsvcInCFzDYrZTkVnemSKJBfp1lxjQfK6IaBOjGfGX1n2NR6SWyr+YCYLQdoFVDhnZawio07i
+nAP9SIgj/TGvvvjQ+vcQSUvjibErHC4Dg6LYtXc7/rso0SVgDGSl1HrnUzCqWJOxtgzpiE/ROth
TrgswdS2oMfdTYZxTBqG3PIEjYSTitk5CB+FKTCsNbE4F98ZX+mePfkHmC+LPBYiHVwCFp5JUUy5
pBncACCn1E0uqD/c8R4GHEXddVrmuR5AeCKZHiN4Kfo91KzWRFk7kz+9lobsxQayvMOZKko/WrUu
uLFZSJVyqTnms0ioXQBNfKVzsGeLsVpfK49PIqqS541NKbbm2oO1LiV4zpiOm4ouMvuVHmi0Z+xp
8dZiOyU+Lkon/CqUEiWgg09fm/jMbiDy+gGAbXYRS63fuMWWRKE25lYDIzHhrQCWbVvJ6FOYVi3M
M4i04YYtF5sWQB6Xx3bFcqvzBzHxEB8+ofNNeKytRf/1jWkdBwdsjR13SvmBOp7s2E1dZYDvq4fk
7oWGGXkyuOXeBzVWWHX8GaUgXRQgLlY/v6f22F7IlrUlcW1TWSa1A3eaC9FiVaqQyMDgFrgaD4IE
mEzD8mRbwFU8BzuNs26a8kTQn2JVv/8XQVd+JSciSUVeBZzaSy1LHEamfNXFxpiAYzfEqXikEE9f
KAglUJctpB7HA3nDjPTbfxTuUgp10Iglg+v0z3kfWbm5vzkKP5XuWW2E/1YL2L9gebJ1qwDekRDd
biyl1U2WTgFC2VqXLGWxoM13ec3uz0H4+vn4s6EbLKhzFRjnFWBO1b23fqVGGCBiR4layfNmZEy7
1c00wNmPH9875IqOyaAv2pyoJCcwOiLljscaXgVUiS5Los4E5/iHvKLg9O4K6rIoPEm7Vm1pivN+
/Jvv7k6V9KbQ9R9wP5oU0BQ94uR+yB+k2ucKoJNJGZgHAY/cZDrS90AHruHAm4bTApba40tzsRUc
xdgz8DjoOfLmSQFDkAJtWdoULLjxJx+NevsbTQmnPQ18BeFkaN8dgmIq/SqO+pePPY72AYmKihct
THSUlQ/NsJrFn9WQgmrp0DzXRLdt7OfGdf4G4jOvdD1lTl2zLNvnACxxx619NCVUiQbG/8YvuTwg
689o9S9hFZ0yvTxnYkc6k1tR4AJQrPeQ9XlFQSzrza6UYdkxaRZmQYugLTJqdsaWPTIxTXwAPXb3
WOkbTNFXl8pjNTi7+sMJuVm3ML19jt2sa5Cg5W433mGC5OWLa/x4KGjaotTdEd6mz5LijUolv5YM
kaINtHZl2c3wbJZojbSLtMHGg5Lt+6Pc/YswE0ZZ/ODNM8m5r78/Vxai+uAdIPY3vrJGLLMHdBWX
ayJ6oC4cKPZazu/lTf55kCpbZavwIuGg8iir6+Adehy0lU8hMAlDm+xgB61ox2up0biVzwyYe9V9
hYLPov6GEpPugdcI34XR1zRcUnaIm0Z5kIOps2j99LQ6Bw16T10WOuw3RldzjJyJ8a7drUMfMLp2
TCOWnjXiT8+RKvDv72gwx66R+TPpwoiBX3Fhs9vfaMshtjSg7DTdtWPQnl0+Y3FUNSH2ZgbQz6YQ
9YFUFa6S6istpFdWfakjT8G36u05gPXRHxkVnDJu99ApqtvIVHFTzlK76q3AAsi9mfmY1Ufce//7
SlQ5IBETzL1Wuhj6R1evmnHmbhBje+hlHh2EiYXY0vM6TIHREN7rtSfJywIyobCIAiiZKBk4w8Id
1H7gbPV4kYPeoL9K/BTfWfSqFxwO7G9IIH/iooPhWgHbbDVp445TRJ9Qs41a8WTw7bNMQc1nLM2s
Rf7oJq4TO79W+n/SUH73qi6SV0Ve2XWhyd6Ey3nNPYJCEQBTtQMm6KkzztpiaC8dJGERIo1UvK8n
DpBggwfFMhOxqXfrTcrmvcuuEbZncKlLxO5vJPZfCaipkc9uOaGJFjbTqHTtZ8LLKEdVYaxqGGTq
eR8s/6nPqz7BVSejMws+D5/HX/iSGkrVSb+VkvXukSIwYVOKOgvbF9FfFbWkNrv/E9/0aMWxmvzv
brvPCj1DyVWCAoq+XgXQM6pAw9XP9nNMdbm+Dn8DKCB+21ChKYWALh6VGeTNCRXwDNc1CU79xQdC
hbKswDax7yqAvdD8KUJcZMCeUHF4rt0OAVrimL3DqfUWarkGgnADpQUP7ouTopXwZttKX4jXssxV
n8n2k7S4y71gS5PgTxb5Py5ALSy/Jiv2aum/cgyTY4Iu4HrGkjbphDzQIiNQsorQ0PEqOrLWxZKh
XU9Bne3EK1G/1/fny5HFBhItjTyKQbSiuViL/uIPyt3f3SMFqNwTtd37BFQZnalYXnAK26drKAci
2ObpCH9Tjji4k6GfcMtQ/Vk4U7Dxcz9b+vspff4hl/vFOCPFpsSO7Kq2SLE7Shg8igcuOnSseT3K
5jl/VF/oEoqYMq54swOTxi5HguJBPoHU/jGa56B6JSzRR6wJa9TXfvd+SmBNxiHVx5dlmup3rA3I
Me/tHV4DOnhbQjHLcPi0LhR1SBBNghTVLgOEHQhKLrMYT+9R1YqBfpybv69BXW3euGQNUbiQ3auX
AsHkKK4Dz8NDjCEXQ565cNif/lBSLAr7/56XgvhlsKsZBcEayzSeqp+KnYgqTJZEoCDrQTYoHIfC
+5+BRZ4esuKYpTu40u78kPCPzcRlqXWnWNTUSxa4Uf2HR03YPgWtZEwrA+/p7AXg+/l28VU2kjdy
B99zyo3cwtbqcdct8nVI9D1LRxU+zMqlJ5TB0i8k7HRKHMTYAfgFsscOmxWidsKhNgQp8/89woDw
XAFa65wUetEZYn37k/Va+nsyi4REsCkR/ftCOuYTLxCR85bu46BMUwXuoxIdDaKyrd37Y9i3Y0wq
0tIRe3zvumROUBZz3VK0rabgKjKRyY/LvkIyvBslsEXQYqGXEUdwPnpafRfPETKSSNEXBQ5Cgv80
MbrWxyxu7fX9olTlMaTxz6kmTKP1x7F8F8mfqOGPiLONog9KIaHykqYXViSFIRRoR+xt4ylCSoBL
MsPn3pawCo1rts3Hlam3HzEjpWQvYfbLsen/FrBp83UzF2BCU/VhNFiapYhZbWIp75hRdfnQRXX0
wuxKEbXPOhIGo2rNqf3CQaMIdop8hxaDkXjSS/uey8YfJllwsoxRPZnBHvS5rb5ih8Z3XHZvfqrr
cLdujahs/BAwZTq3r60IPBGKb0omWA3TfmsAwAfhJx+tb5Ha30zoGncIqv4TX/VcvwOu7VjEk1qJ
0EsZmpixMnOuAtauWPgQs1VZPS48EQCgoSkst9oarNC/EHA7ck0cMt1KgLbUjtQ6yUYVazF26cSe
02613ls8eeVcpfWU0Sn7IO7WAB/XPJodRAd0Qh3xBtNKHQGWY+oUOW2h41WG29rwfoggVX+pPjjm
2GSUdxJffx1Gpo32dgw3L7Ahh7aaVSf+Lzz7eHNfzAEgVrUZZrWAy9//mW0LOJgKxG0kB9I9ZN9Y
jAxYLrpUfr8ZXUnTtrlTfpmLHQ7xYz5t8Bt/KxYuLY3WBoXfxVWCGZ43OQ667FHBHTryOR9hUkIP
bcXLQG3tNXXtLPKGdV/K1ISpZc4B/zXHM21ieL5fWEyHcz7+J/+USo4aSILyHR5k0mGf8Nux5Lco
FPI7ZxjFhdBS3JRxRdQ382VCmL2dq2PE8iZ6W9f60KPNAFX32xWsta5gebCgytSGbIliNSLW3Ita
2Xr+fkITMKz/c0MHipxjvXqTgvRVrgi4lLZV4mD6lIOLUsI3mloqxwpZM9fdrXU/qyXAOtKQtKRo
4YU5MQkV+TZI2MOkopvGDe6j2jD8siVoqljJKfA9ePvxlBOzk55v/iI/R0u1C+gyYM6vVNoTMiF1
A+ZOWDnEpesVAzXSnl1p3DFObpBcZ9hnhypDcMhI6JJJjyk9OqvdDJOLYCOCSgI0NjlZ/TTK+Etw
7T4AYCzirULo4HkHVxYJUbWojaIu+emrEwsa9ByXAXUui0ZzCZ0sZ3nLx4CQOO0LDtgtHbz1Kdya
Dbspgmg+ogl6uVQouRrP4fYdRyeEBaQAASZfEDdUXGigIGzn8Ib5XtAQF4tv6jZMKUWucRq5r2uf
iA5sSZxQdaEfqMZxVNfUc11HOcZZWh/2wRhEjoBgWYRvJZvINVY3AXOpbNJ8lY3nK0GbAFzuQZZQ
CBz6QiNnX9OO9zM2LMxEQflfbXjHegkLaZWGbblKTK6caREMZCGTwHDg9nnDDiwQqCXDE2HIuOxU
mI5RF3lF5X0x2X1h66zVR8Tg+5oK2yrSyjAWB0f3/h4mYDXSX6ri41Fd4Bf9TmVvbbkmMLBfPpH+
nSfRwnunE0/WTCmh8tewm5vYklYit4JbjE359j5kpTd+g0q/IF470XxHGRWybpzhKU0MpiqwgImd
4HZOky8sX+9UlUiP7mvzT/DrTjd8+phwOH4G/NsTIb82R3AE45IVbOH8Vz10UEI1fmEbD6vuDHUx
S2YOMExvNzwdkE06cJNpjac2pPPvZd0FX0SdoZoVKZ0nuWVZ9gW7hKFWo6/XVomJh8+7z/Jq2H/H
6mlbGXNOD20pmdaozKTcSI5mUJM6knOK+2KfDdMeoVGJKCwciglQttiK/YkT4nMogvXfXT93Kq20
oAhBP4xi8pUD6fJPdBm2BegTPwoF3U5apGryAShaPahqQs2KkEIGes5WKbbVHFmU7U+F2bbKe/jc
/LemmupE/dWsxVKHbglJCpiNDFwtuoH5PTaZT4LUBBkefOs1FffoRz3k5DFRxeUuYlby6zNfFlBc
IRuYc+0Hh4Vwd2976Kf8x4ODDg4nT38JhP2kEp0ZbAsLGWfUxx25pg4JJxsg1nY+EDEUJjiLWtaU
v48XeEgroNTe0O6P9Xd2DEGNW+IqgOeEBEDUZYvTe+MIlhTV+RSTYd4Hqn9p3dGe8iyVP8So4wyQ
p9I+olo21gJgoXJsJKayJDkZgl37fCdiy+ntFMEU5ha0z2AU7MdbRfIyQQd608NZ/LncB9wNOy5H
yMvwvdO5SzZPiSvDFhwJk+fZV4OSJY4NiBtI3zrYS/zNN40vj3gNCgCpeeYyKJQyOeRq7sYWqt26
GDbjTprI2Zq8mwrOhwncGBNNh/beIzQwBHtbTBWNVdC0W/eQWgYqyoBKoXWfemwG+t32mtfxIXRj
s8SBGNehw6PfLb5BevP4TLiHUl47mNPItcPcWUpy876oCyywJYvq/U3K1seYRsvXRMyp++MSLU0J
OXMZJPVVkAWAGLTD6gRD2QLkzvM7AQxi5HzmoQdUOFsEIa3z14iyYpxEMAztcfMbPrJ7rey47DVy
Npq4Dnssm2JVuMasQYxSWhheb5lJL4Ju9n/K/I3U2AhglFPITntqgTlHLiI2td3V/a1Exzr1oXTt
66hMqkrZUiy4gSQ3AGKJ5c2AXeV7+ux/9UyM7rNEkvSaBBm2mzijYg9bn+Gpt1CQth0dqWvAtH8H
lyaiCueA2Lw3JWJ3/2hsjI21B6Ki++FGoeVFQs7359422bLISd+7SHWOpfCyHadRxbfec07W7i6M
nfqMrj2ffPs6CeHBfbH8isIEMYEFxsdk3AexQTZBj08qGRNkIoRa1FcWleqf5dXEYMuHhjxEkJVC
l4VxNjfpSpWVjJCocL35okAZRRsCaL1y5qY45WRBYi1LNblIxbBTdN5uhSO1nNBmqoalAtz4/DBY
ltFegyqNemlkFkplEYbqze/ufiUHw40aeph11BKC+Vf6l6YxukiwLVUxH6HtgAyNw1wwKvGN8C6v
h388r6fb/i6Jy/pkACmIMpGzILB3GQzQN1Yix8DQU5Y1ggzl84HOKPlVPUGX5Ji8QSWpO1lX2j8X
9Qz2/yKZTR1bqkWiefyzcbJXdll7FqZGtxKYgQGK1u6MPJBG9GJ+5c74z0hrpJy5aY3oGBLFhas0
r65/M9SJ1rHBGufjQb3Or9rFkU91tpvNGWKwqimP2b70Q0eSMVEa+hsWZ34CrDcIT2a18FxpD2du
qjpoE5v7YKJy+Hn6j6e2dAiao8Gn6zRhmNECWeXI0JJ4GURufpNGfNzH0o87/yXpn3LhJC154NbJ
8/gIRAWRnNFq+oFMHXUDHE2hA5pJargCw5Tdt6nldscMWOCTihf/kUsTCLOtq8GP5bkYs7/aF+cY
IMeMwNNq9G1oMt+8RQ2mnvPwLUN9rAcAuYApO61OAACXxqrxHo0IynRT/E34IOUq8U46q2RHy4Zs
bjNSol3W3fPbJJd5IE4TFocm10hfsrNdNE98tJmtphEclB3MrDejJhTfXijLtNYRiqhPzGH5poqI
Uh31Jjr0/v+ufHKw+zjj8oBdMNDntQtH0JvrIK3eVEQSqIR70iEN2M0pyMER+C1h555XN4lwFcXx
fpDx2nulGVQnt+BmKW3yFra7JkH20Xa5vU4c4OujwZrElR+z31IQnmaTZK6Cmfn7eFqgjrpK+Bdw
crwpAajpANRPfw/s7Dvmr+zvdY0v25iFkAjmvUtDeaO/N18QAJ849RHa/cUhPcM9pzYbDu91QZXz
Nn8sDaioQkdczx+0kaX3DvFSBGZbx91BX1NavSOzk+6pVRTnbpLZd3XIKR5EZ9zgeaf0xfy64nbT
3Np6YGmuCfxH/Lr/MBQPY8y2OYRahKBBc2dN0p6bwvPO1X+zsqyYO9l+/FpcZXtmsbQ/KrwXQhv4
MmPzB0qITfMDSNOhsW15JGWOLZTc0rEBzohUUutQigdl73uomc2y3lmmVibJl43wkSTR117J82WZ
cJl4f7Joo8ulm9PyrAzgaeW2GdkZ1RqkR8pc4dUl43xWHXVfYvw1zWtmgUBPPMhKSmXjgGoEWIpH
z0n5L6WCzlNOp/q7Dqc5Dya7kJKtSb6rQS7sU6PeXPL/hR1XHzlS4/A/c915ppBVoDy3mScuLtzH
/jqZnMSUUYijolzvcFjig9wBJVjvM+4LdzCnQ4oK5QJc6OQG22Ys0NtEdj2WDZIYfdHYred2SJeP
tBuPIFQ1BYDSsgdRi+olo5LAbK1BHT4UQMUQQtI2+PTAuZk//yVzVHoHqve8Mwa1qWS1YNNx6heI
6Db5MSpP3bBUNt4C1M517WsASIY3KOHhRNUWUEqTDHgqG7+fJNBrijBP5kmKuwSeN7al/PABsX/i
YEDvf6HZHf6pCoBnOP1V1J9wUGed8tMcWZ9TzfS04ehcc2ycWJdcwl6dl6M0YsXk3Dw9sHBVogi4
DeVJWNwZkDuv+xxjOYuYexhaGVwwNfdUkEaiZUtsr44lVSdUGzxlIjdhJeIlj0A5hR2TuPC3FV+/
w5ACirjFOMdvBe+qGrsRgUtYkRpG6sK87dLkBz4yx75jwVGghSvJnT2gtqc4GXKIcHxclrRWeUfn
prZ1nPng7/oW3mxg6BRgNarNlKysyGZhwgGsAF6cTkyPAZ1372L0MnlphKVz/7cFg5eq3NT1HJUy
zFGkfTNJOhz4y4ftInsjhdCV9hYdp+z6Re3WEv+viA8o2ivuufJJsm8EoThzFCoivdU0i5qf4QRH
tRv4sf+T2Ce7ZW+S/fULBG1yXQsJLUdeQeuKF8jdFu2P0SXgf/Jg4WzGR/6zNhgGFERaROfzBzzf
CpGsU2vFMpS6mRwU0nmAcwB37ax1KWtRr3jh2ZkaF41OcysqPuDQeNa+ZVDp4/3vjt09mIBfcJHQ
WdsNhE8cQPC49XXolZX49I3fcw3SBKL9mwEDuvulOp4mUQVdYXG1rIPwPYrRnGdIY0awiwFe4NsF
sRujlS/XzwmqzczSoBR8X0MC246GsguSHQglfxoL9lruuNosYSO75gq9XRAmdgJol5czwOWs6kQV
HRsf79XAdA6BgWPkrFh3fSulCKU6UI5d0pSXdx6QA3khY1GZTSi5sABh55rcG9CD//NuqMDUhoQc
3dldgk66sYG9sglOTO4K80GgCD3V0x7Bpq3aV18YlEu3TibrMTWhxlxExN2r2uZwtYuztmMGxMAl
JN1P06jZMGj1eEPfdELwXOPkplny6qUggsXMfas2ihls9FW3u8sGUW/zIYsY6QRhgub2yfc2Kz1l
SlCdahII8ItCyBPwTc1eDSRqH+KbZRvbiahoicGcTj0QusRN3i7IyI6/nNlKDUoTlP00SYCTofMk
X7T7n4lnfzwHJJh+5D2/LuIyON6EUOAirZTDcvAYcHPVLKujURqDWFndZqME8a/QRnnJJtEAASAl
Zj8X8MuLWYQ+6c8rm7x4CCahhW1BU/ERnUCS8kf0bTWzx6HusSO2aYF0liRGl7CxKUZOqEpatj/k
Ae1UZkablhZXkN9x7AmL1IPiXBCC258vVlm/TmXBG0NllwNbpDOH4PaYjU87j8BQxlBvNkXW8kVW
qDklBj3R1RYzWB3dgIdhhzU+3geNpBDxRHzV387DaH8P2SF+GYeqDH7zjqHzEWQOjweygqwjw6jT
kLQpZbVdHzYchbb1CcOegyqdDG5XnZ+VpKgwrcx0pRoIMGvCn3D/j1hO1utT2Zcmw4AouWS3A8t3
vPQLlCuOOnxskZCgaNsrYBqEmHZ6Dk09RQYOAsBxEV9qKAXnOf4iNhg8nX4ARegPlZmgq9C4yAlS
v5gYgEoMmjdUHK9iVjOlVqxnfnLdnKUNjtwYMhKLeNY2lIVCjUd1v7Yr55HhFeyPngx3fkpIKQJs
hj9dE21Q649+sPaCph9iRUhKFX5W06nv+Z3n40M7R7HDdlZ3u+50q1SZo1Kr5fhinmUWRLSMZvhQ
DX1q34E9sbSihKgpUJgkUCF7CJ/7H8um634u4EyU8pX69ZHnepu6/h01dsUH97/gcDuPymWu2ip5
17SKcRQ/TCChnv7GllP/2ACg1dz7VmxqrzOR1YtjNvbTHT7Gfi0C120OGY4ZNYcRYz3qpZbHQnZK
BRkTWv499ZtxsvwRSeua12p998vsf6lWroxUVyIGhwdHsvHAujqp7UyfbYv2GqheAuTK8Aik0Dlk
Kbfx739wkqP+Cn+2AfUPvGVVc1OBscwhLbzwTnETTrjgxnR3Luu5oTGDkdKzc/NxU0zgSizf/PSl
boNz89PWis34hroVNt4O/06jcn2GFRZcXYSFrZ9AXfng4anRy37juWycYkAbQQrWlZj6xc+vyMGw
mlZwDbgKitciPL0zIHJze4VoLXJd4TUxXzB8YRsDjfVT0Y5F9+VWxLtPV+DeEQBPlc76GWK9mN0H
OpkK6Cu3+BOiSY2IhpN/WirFFyge5DjxLAPQv5uMIw4oHCBkdmIqEbd+nlN+URsc/lbLb03c0N2u
QVLeuDuwfP7a80jhpxoaj78dKEMNKUQsaPSxOyNkZn57Y2rFuKqzbFUgGdgvDRMjgJRbU7FMWGdB
PIPiZ2JuetOl4yRRCSLi7/xJzXKYwaRM5swHB4aD+8EPvmLWq1arZSp6cT2QlZtt3x9cbpcixJn3
g05kSK8PG1VuJ4ofa2hHGzQ8ANvAHXLGsHUEVm8VnluAuP3QwBWWHjfxZKXrJ5b4z144U/PTI6MK
BPq68fDiA54gKH8lgHYtMk+wvGn+/nt3q56ffBNModIlnfrdVdHfbAsPs+aWKxQRPoK6RPuxg9cT
eTuKtMS0OPN6muSVJfR6pL+e8/giJws21LCKwUIyG3tUQH0wwjQLOBo9GRZKhlCDnhIVwu1QjWi5
gdsRVMNFDpYg+Km6/R218P6d/hqqLjpr1/N1w25N3XizUMFtASO2LdoXPOeduB9s9Pv5kKDyM9+m
pQdGXG01R9AaxQhTAPngIN3vFvfn+coVXkNL25xpTU9LxnU1OYu2HMPGnwewrWXfFHN0i9H8Nv5J
zafJip1l6qS4rBJHxTO40oedw6RnYlu5nAaT5+mCK71e4/vHtq/ZdkwHpfo0QfoE224GVwourMgi
J4tpwSUXUfiWr3YEbTzRcEKFqu1E3GWOCEaqYpUzd0RiWMzKNQuPuGRSh9khVNkY8RWCn3XGL9vt
+ioJMzIf4vQGl8tuaCKkaTkYiRWE7fyKnHjTDJr8tFhEkSxJENWQYpQZEiZQwkBjQm88je3byM6f
BALmK8LQcQD+P3SMetr4mkf2r9oI4SUoAj5J4kRyG2mcP7BBYMTm4QUr0I9hfv4p1fD0wdsDx+BP
cQX0OwFX1of20ETKvYfzKtrP4uW9/tCw7Vqbhpl+rnZe0SN3hD5HY82YRRynTRkUsdGLNh7Vx8pe
g6GaIrfP53B8WAEX0DKKTwGX0aFDpUFhG34aocls3askvGiqCmzXO4ZqyewyMwb1SzWlDiUZC5sB
pav6XBWUmvTUOP/QvQNldGGpiYkp6+9/8J3HwBrSMjtMzbTfW4vRiUvYi4S7PyThwm5/UyHBWn+l
zZGZZSPwVVJNlzxWY2I4WfcQeljSjJFi8lRovVzL6QV7hQ40UkjypXXJ6YuEb5508EW2yg5sXpnC
nl8d+4/fwuLELkTYk9DWqR9wt56aqakCxCNBYGujQ2nmv1S0kQjUoc/qxk4o3jMoa77lE4275tXj
XsrDLOaNhqV29r/sMkIw8GNi27ToHQ9tzqZDhqwMIOHlDuQcIhzNud5rTgWBufBEtK4oiDWDI3aq
K9N9APzqntEj7AzX06wnCe6Yqbq0uyEqdbci1bEq0y0GygGcAEqbDTxfnsLAIsIa4nr9OKmjLpkU
NyZgHS2K7alsFRAY7NiUoYpPTTPHkETj7J2q6yzhbIS9J43MSqtFXFj6UlLl0PI6x7krHoP86806
yu9m6o1+tpqm4+qd1KhArbXNtGa8+An4DBLXJdUBsNBadw75BIgNH4QK9vMZ8QEGQNAUAdX3EhY5
b0gTXteXuIjCchE0K7yMWJPtApn3iQOCzH4k4IUk5zP6fKd4p+yE3je2iryb/j1mF9KDFG5KC4iZ
g+HGEPfs8dfx41FMuIihAlt0dFgYFzyUMkFXkn6MYk9P/YD1mS9/3IfAmTNLCg2Kdc6gN75Z3RmN
0jTrmY9JcqiXnDV++gB7rXTRkCwd35SrbafHXjg6mKZYOF06RkHstVJF+7i6wv+hf/gt5OKXx2kO
YLtgOTBhlYfuVVR2cC2oiyyQoGJ5Tc9PMsAz4lape5SLlLU/CRCFtQaSdtIf6x+7xnYXY4Mb7Z2r
pMhgibl1XJlKdCktDSlzdEbheFKnpZdxa04b+2ApDX5/0Kq6M1dMP0hRS/p/GL49uS/T6y2tHl5h
TeKH24Pwc97SYJ0xCFwn9WCPoUKaYsp9DTFzfsh+crvFgLG89I1CXZ9+UVFqZPg3CWOJk+uf6DZb
FPKgqReBvFJ/uHbhpivAmtO/A7smOsZzUoTxqFPLO3YSLy+znqgQYomlZN03QZpph77UnImSp7qf
azIPJWw6I+jSzKaVQDZH+oam596k/SceTI/7z361+Gl0Pd678OsCB58kIEqLXmCoXROWbwbQK29p
JBrpLC5tjL5+eY8INBKwZyUu6ugGoqtBPxIH9cITPFsxmxFQBN5cIETgcl2MICL5ARLiZ6Gzmh43
ytNyEN50JFhNWoj6VzhuIfbseAqtQga0MMeJQqq8qY/c2j2Z9oD6YMp6bGDvKX5OLnGUwf4n05wb
MReCFYsvecFuU+iHjMsWJHt23oHjgoUHmN22aYo0aPEAsGrebyPvVSOWMoqfT/T8wrTXrqnHflGV
CiRafPLODcLyAfAj1I0Rnbm6h/HjIy6KCiqu7HeGoiZMcsp1KWaSpfJUoq/A7Ge7qFpe4SuiR/mV
06RbkU5fwpNovjAohjJxs1D/OTTXjYsJYjYsh3k/LnJH+A91vMNTz62haHmVFSucTn28yM9x4LdR
cbW6YEkz9QTZsC7BSZNy9jRBT5P0PKCgv19UpKPJdrKvtuVkP6t9PT/kxs9BkttKWspW7oTat6iW
8tre5XU4kJBDLtTxMKFUO4s5OJqICJduDZgjld/OsAQQhOZgXUlvQ3QfhurfG9FNVeftRUb/7ups
dvptVYqYghcEcSh8P1V/cu9/zfWC3de7x6xJzEVfO3KfCPJH8l3ih/PSD0g2ACeZEfhHwD4+1hJF
n047PkOau/SOr5A57W4Ovd8dWM7RiWLOS7g94/1ok79nq4AgSTdMCaXxHrF3KdXnwHbddNi4Ziww
eCRIbBvYrK+OlZk5w+pU9QTTnjvWnUXdtm0NfSClgf3YKPjolzgGhw4PPZt0mkqopTLZscrksSxz
Bp5knBDWdYOAade1AQjKVI0X05MTKz+yi2HfG12UB3AvCRxBLbDRjSly1Z+GXtmClul8hTzCMRnR
Wc789hVhzx848lqvHD3qmFf+pw/9NTbDKMiULpgyGrMmxFHaXykjOUVTBqR+cepwCTPAtwickQHn
Xtxsyt1oDQxtXuN7iVFJndLEbUKTTVR03mMjaneztNILQi6tu3qO37ZsPlUMyybmvqeo/QJDuOyN
BO/nbBADCkk/o5S9YpXvUUYjHN4vvOGVvC65fiQbVtxpksJ1DLSBOapQ5kHk2aYH6wD1yG2jx0Gm
W9emIsgKvDK135aPd8W1AOkCnFn4k0L8WuMYDFTuOmwld87oV6EwOyKL3+fu5OI9wm92Ec7oDFwA
b+L+ZiqewWue1Vzd4PAswVFcBr+7TUqAbklQCQ1oYBKs+koiZ7r9jFn8d8pJwIgGUH9nB5o6l8HT
DZMYuaf5tnHxE/ULltstC4SaFcLqCcb59BPELWGmlO3emmw+VjuhQ++5KHCT354nee1nzLS15LVQ
XiKB4dLFeFcn9cAEcKLDCY2tQx43fqewHOCZ87WHTQxfIYWaUDbXeAhGgoFJsVVW3la/zL4uBu20
pxJp14PC2LEr9pU2nKtrb6/1Vba5G42cb22VM4zhECMV1wPwiKO+lWjwYeq+FnObyELwOV/5TZjt
+JE6zdRo8BZl2Mwg4TvLde4oSdzs5SmoNX4JIQBgvkZKiWMVGWzIr45z7E3vARMBMpp6ldaIFVhd
TNW3/yivsu9l0vVpZw2VCT0dGrqf8hnhAruVgorVMeIeKXj/aNfMKrcdnHv1tDnnsFGCCdSI7igM
0mP8ZIK4qIIBN9g50XKDBp5hUjOkO0U6GVnKljTLWe2eTPc81iggdfiqbaAKV5N//XLp5j/dixJl
xXxCE9aBZr7bRybDC0A3E40psZcD6+11f4/QFSnKDiksz//CzMKYASOmjZh1/zMchhRK/z1Eebkh
HT3g9cJz8zhqBCChJ4kTezpSNKpxoZv5AL0EJPq01nzzuD7y3kuARQjrU+Fz63NNRVJjJCsUF086
JBaoQqkWKTo3Nr22XbGfQAPNi4dvdEkHCedsH4u5emjWqjL+gwnRIjywk9g8lRKMxp7gZAmavyOf
pzUi1ClRMnd2FALb/Z6eTjYReAniuEDOEwjNMjh0tCa/1WoH0VT/4jNT4C7gOuiFpnvCCw+Boyhs
WibL87fE3R9MN057lSFRbOUmXJXivxuntOzJ4Z26c26GsUPgb5usNNQTCcIM44A44EDKkhTRmwmV
77HMIlwHRzOlo+2TaGH+Wm42t+ZhrdkkFRLI7n3T0toelKjp4xT/WBlny+JjS4AjCKqvfm9s1bCk
mDPBvlWoPkEzNwvEduJgRPqVYWOqNap1iRH3wYJ2xJZkjz6j+Y0DIQaifBa+1PjFL8gSuZmi2KWY
G3uY3y5nyY4AiFjVBm3g3fmkVqc+n9XmnawRy3H5C/EbXDc/XVsO0EZGNyRQSbejlvbT/TEKzkv1
ku2qDqO+1dte0NGO7wB3SrK67rUX8jPyYhbsjyV1OcuKDcX7IvQEfoSr3EogL1B9X2iUf90/jRfF
weIxzw45DxHlRQd7K4nSYXI4YRUk5BM/KfvMMhNJeH5/pUycAtkMEbAIknbsttmBckeDmvu9Az0m
gK61qmuo5VfWNQbnLNM6mELiLpMtEqyiUOxrhmZjoffxIkILvwuoCDeRkrGbT+QwpuV4sEpE3ZD0
5P8ZOuI12juaMSXgJ+b7LRH7cdOItQ/8X9wRoBLz0VsckKBeD0BlMHe3Ui0em898jDEuOKDOrM29
UQjqi8gelyXkvQ3RSFjBu37RPGDqD9yfv13xopjxAl8U24ofwxI3yNQMUSa55tNLxrhok9drJtIv
EEBUbuboitzRL5bVpANQ7OdACNir3RtkhS+k9a7J5t7uUIx/JTH6gMXuejhOiPfqNea5C2Ra3eRD
8zJEMDLnWFIKo2Lic4toMMbmIgfpZeA3JyR10UskEjZ8ZFEfIjANxCwpsdTn9s12Kz6JSzkECOPj
P7hmgGhCNmH0qoeedwOf2/dDqV+ydjMyMri0wu6S79hxzmyOVVdIrVw6a82xBbueAvHOLAbC/SNQ
voZhbiQQrU8MjZQGPxdTef4b96Oy+3ISv4nfEkHNVT5iz83CwJQjsuYM2RChftzNyc0Pm/6SeCyo
m9DUndNORUKvoU55kjC7noEhtxj6VX3y3gfGX5PctTIgJSvceRiaLubvxjoD0/QqSf0dPGKc1uHw
e4g1HWrhAykh3xEcdzYuhb1USr9lBb6l8c/kfpcCnzBbVwuh0hT3MC2vnndrq2Oq0B3ebqFCBbnJ
xC8e2WRjIx6jWkuyrrNcDyRPa+uBQ89AWYOkIJpD8oR/PBzDGHv5MNdWzpQl+oXzCs/m5hqcKZ8B
0CnNdG7ZeQ+AVkAZh6vHsTqpBeGkQkQ67knoM0cGXku9/gP1uZUaBAnC7gI38QoldC0I1Kb/cAbD
AbrqFfI1VlltHQuAMaNorSof/28tJz3/EHKfZYvlrABjt64DbefF2hIUnP3B7ekPI9lkiIoeV2iU
oujQHBhwOv5P1HU9N1gYjk7t2kaLYXhn4lygXOjFgma5bitD+AnqVtMmaNYSBu3IyesHpDeU/qH2
gBIDwRdQ8xnFLLbH/SjS6sJGAJNkHwnsOdNiAahludNGekBroe/guezNA9qgJKXNvpu1FO2yzUYs
zsx4Ux204PO5dYgpRgBZh9wedoIrHS86FF9nhiSK7pMCkGelUCle2dMCx9y9qrwLP9vY8n2rlYtZ
wFavy7YNpRjBvDGZq8P6AEGtKVkuYMJB/kBRJ6JFBxErPBiQYWcBtAGqN3sGxrbIqWvPW0dOS4mz
dMT3cV4LG36SLRw3diglCNv3MoPHdZJ2Mc7k7/FAcWuow1rBtO4Lxx2/j6/+iu7GbqAsktjiExQo
TgFzTOcpry5CYaialJcuh71F1C5/nkiidjLmVI9abu/5kpqDWDWdw+7kfXQOmiPSNKir7UDLjIaI
nTlRwpzIwkZeh7y+SyQNDDSRc94m83EFLKTvWrjnJvLUfhQVqjCeEvzwAPhmNxgNjSzAyYBVkp5X
+F1n6d/0NxEivCqJpswa6Q5vHO1WIFWte8iuRf6yEPcorZBWuKCR4rRs8c0p2zipGN1Z3J180xSD
GG40gcT0Q7ts9JrTzIhnSlrn83iilnLMJL0yh49irj7IYWVT8dAtXzvBj6Yk9Dz4AnOTjkWzDZ2l
+Zl2TDe11WDJQFwH6c9oqttezKS5OjyuK40dSAg5djRIyv+MTlwB+SiX4STpQr/z8YHGVO27hwK4
UloNIbtfR20JvWAlt0GWQCBudKCK59y4F/h2KGcoVPzwy/26DkQpWaiIBPsMoMJleTIbNHOxpLg1
0O+cV6RlzpkAr6RqepZOUBjKV6voUyoH7l3rYJQNcnHi4l2euXDsmPLWE/JDvdGrXSRTtGOcyz0t
Ldm/6ffMosyuzmn+fstI1o95U9/wzeNWLrMVF9nKsl+wJWSdl99lZmtgQlWGKBdZJ6/6cFE3QV02
x1PPyZLV0bMapW/uSpeW6R6g5y5/MhZ07UlzLRr8WYYYF2OihA8q8f8GOy8mBpjR2opV5RIp/hYt
YFWEvTLYhslHwiVaObupWq8Em8p8H6C5Hbp8GkW1MX6DEQX84AEO4KQ225XvGusOxuFomNsbQS29
udETsWHdNUaWlT/h3dlLe/6WFItV5jAtAkBceR0tt5ohkavJwgD9/UxZ99Gk+tK9hG2XfsQY+DAi
g3sKSKdDw8DtwMXARNygsUbJaYM29F0wVGaklmf3u52IQkZxBWIbQ3IzbZEIblA+EvK5FA55WXwb
vHM2Dk5rR5pa/rmbnP1jXz08twZh+AQJTbZJILnVN7NKy8gCAA7E9Sxk1ELpBIsKtYZIbUIN7M1G
itvOLfJGXwHiidBwWTJOMJsdqamvw6S2JxBr9IE3KJEdrGTvPni0yS9lSbEx2zS+up5rnu7Y1UlG
PaWlkcGoku3pQ6dLSLclyB1PbyqmUPQ3q6K1yYD5L3yUXg8N4pa7jYG3fV0Y112fsZsKirZP5NNH
vlKpKR0Kri+AZScm6PX2tjI5HVp9GqIZDoPs5lAiUa+z9v6LwE0laS0O7kqKSANdthyYSXps3K2J
49B4Y3wMF9oNoqV3fsxwoGO6tBxxRTKFcqaEDTcCtUnNp+yaGhErLsQTcxXcRm1iLYzL9jgE0Zra
HBFg9cH7J47y2kt1OV1wHKKS2n1bMtKKkrlsKCJBocqMZZD35KLmHb7/ubv7sK8EhqTX9/NpxlWr
QcTMEPwDckhGWdPn59niiWGuDKQC9xql7BqBRSyqdzONgVw0Fin8ThEto5NAZm0e+5cpJoIbjWhn
e2DbL85WlkdHflU/sDrNKEJ7JsoxgQ2QmUQV4safyBGwzgplNP83MOmjyxIr1oZQAKHURhfecXt9
SiNIA+dZXmh/a/Mzh8VD5qd7lzBvyM06ZVuVVadi/eVCj5RCTGZ4z0dXN4oSDuVTdfMQchRB3N1g
bC01kK5TOl9f28fNl9JWlIP/oDX4lnQQuuEJMgONjZU4Y/hBIQsmlXahoE81hJrT3g1ElnBsuOsA
gYePUUV5X3cjZm0kZJRFmuVA9PT4vjTJdlVpSe8bD8ybfhWyrJxvSnkbTQjdTEz9Tt1q0iYrnmYT
ykUcR7newZUM0w9CEwI417Izxn3ZSQg1tNy33nfFeWnioI1AzWrHM37k+pJ/LBAlFS4zVlXKkghB
ZQV1/u8a8A/qUl7+8CcT+AFVhlwXu51z4YDNkwIOc3cTsdVWmiQ7GBQ2Rx3Ws0nx0MU9kHrW+uIL
TOl2kiU8mHO7boXXkD19+u5sLw6VilgatpeAOMLQ5tF5gAbMWfItSLZoZQVrwWdHqcEeXUVIDSXq
O/hKRWf3G5tzAqnnfn4bub7Dh6htDCW2MIUPbkd9Ok/qhagd0MNu9hJLAe6qO2alTvF5zXaInMC4
2B/yagLTypmHy6s6cObW0YmE1yFCJMn+Xj1klRzb80M2BKd1GsbEJmHbMoLeKRy6jgL0A5kZGrIr
xIzmtzSNPznawGyaAZz8gQ3o/Cv7U//JLxNGIMWRP5IKROiinPsf2v+o8pgMaEfeI/vDb55AFA0b
gnYmCLI0ppDKI/w8WX7x8h+zmMTksSpO6q3Jn1h18ldA47HX98xz2/Bkb2aA9UypF0L6cea/N43F
X85KbdyBGtKH5c0hyp+m4PJee5vMFTUz5l8NPnA9IOSRGNLWyi7xCPdf8fsBgw+RP1T46jXMqF5p
LfvwPux2wlzmAzFhAJKwAqh9BYLpPaCJEgkJs91Zv09q4rg5V7cwlnYXoZdduPftxfSFUa351aAJ
pLhurnTULiWpvPqG+ed5NvwgStXWx8dG+WlNG7VLR7WgCQuJ9HTuDJoTD+rA+BfTNuF+NOAoZ1Ev
zLIBDVKcuHIGtZrB0pUYKYNlFpJhUH6UUa4z92VGa97CieMdhdP6aeUA/IHa/rsAKlzVI5JaSJDd
DwDJ1FUckooX3JNpXX5+fuFT18xtuBv9xyrdOuunzhMEy2B7rUKUoA1yZwVF0C9ZiJyldAKGlnDT
AB7F66v5qGhKApsQn4YH/FWvzy/9XiUI/AHQBFRryfuZlr9oSjbo3/M9FA/oiLx3jP+0PuHkyNgH
ygWNcdzqnCeqF/YoNyPIx6LR3bxBpB+rqKAkStJgS192Gl9+ceMeylYs9KgxDd/rAFoJM8Vf2LkR
op3V6uzxFJgpbfoItn0FqsHWzYIAoRCLbHTSaMykvS4aGnnKqpOKfVjKbpXrS3Im9sSI7xNikr8P
jBwyvlhSq/ws8mE8UGYOpqLJxGgKcb2Ep9xGB9+ccMhTWI2B/MPiogA3i2/qiEwzRJij6fg7KjFJ
Oxa6VDa+1P1EZhmFOl+y4Ul8KaQCvFp8hUgL5nWMmB0b+IoNQEreuKX2eu0swinIm3Y8VHxL+VSh
QeToGcMv+4rIC4+46gTSjUmsJqxO2FKYJx+BskXYfnBU1JGR079qPQejJKYrmcIpM9RKc2t3Xj8i
FLVWzaudLPajOnUoWgOPpa82MKDCTrOS/nF74y2mPU2JfTVCqgG/sKwVim7oHZxvaEgxnA4ORZZ4
NZCKT6grp2asNcd5Ic8UUtMi1pjs4btN42wzVxrzKvY3Il0hkCd7+LgFH5rT6gVrlvyfbnKffR4u
b4a/HjOs9gY4Dzs2mU/2TAr2ebjfGKhNce+ZjEkLKlliBjQ67d4mDeFr8NTZ6TnTcbOxvDLu0ITe
87gHzR+VuQjRvHQ6LD3+bk/DYB4s+OYkqevglrLUxxwcjrn3CbQrmFdxUu0Dd9EtefTtkCV9p9zV
N9wj8MUjh470BK+7dTLki+PVM2jYoELqY+438tnytFdg9m4aBgGxjazk4/b5FlfbePbvT3KbTqX+
/Cg/Z/Ec47/6lZ0QhYnWHAQHfOjpyowl/+7oBX/zUJYFxxpumLq9PG0AWR7KPJF4Z6dfKe2grhQn
t/nnZzGOV4+HmuiCAviZqSv0oOZpWBTUIFZI+J1aH/xdKMyN8e8Rw0zVJOVC6YEgPcUuGQD85Sy8
0o9TNOQb/yuEWNCN4OsjDwQ/8yH0mNcvwnq3+f1VMulmXwJoUi3kswRAMS2KDfVCX/dSGbIsQTta
AA83IM0+mS5/JJ2DKBFaaWRe4qcuFg0SOOV7CYlr/rutMI56J0ELXyDVa+eH1aH3X/R8Pxrbcui1
ZzASEVcYzpUpLjU/V6MgVELWAIjrmPWyoCYsA6zPQPoEwXeUUj8THgebwaMnXVpM8Y/4KBKow0Ez
opZvcexxOBVGYy9o1fUIqMcAP40WCbcK0zyEJIO//wqEDOI7gx1L3z1WOgYAbVeIGvNDN2D4czqM
tKCcbbHFgJJxaroR61YWvLPXW5DFxTLIpfGgkWan2hUWauGvWzQxRb6y9HFMqr4QJec1sy8S3kaX
9P7ThckBoBlxDESYYH3R9AABNQ8Z18fBjlta0IsxHw1kuj7aQv6I4pktnEmnKn4Gyr9Ep4YB1/9l
qVKvwHYQOoc3tkz+zegS+z8d2Pwu2XGS09bydbNnrHIU8BL5t3Rnqmv+rS4rLN9N9lCeDl30MJok
i7S+jb2AU0aGniT/kQvvg8oZ3gTC34R00H8d5T5cKixEYBhvc1kDWNVQxdqFLnU5iue958+oCW/i
3e+xEKBIjYSzHiKvGN8o4ZagtcaYydMbBE1mcaoTK809PdyG8eQkrK0r5VTDryHGdn9UI8u8u9rN
U2rzV2Mk/xJlwwqxDKbq+9v+dJuynbc5z9qunjgZweNkmjkYqt1sHgRM3e0Rvd5z1iCKZQBXLv0S
niDVvjv8NcJ18Q0X7oIjiqFdes//qpKen1zTc7rtBdOQMiOLDK3k4WmOvpT/DTYEZ0MczVqycDI/
tKI2RnbgIhXH7YCEflDPW7NFIrcbH3fur9Wv+mg8kbkfYIfjkXR9u44PfD5O6fn6i1S61WIsFh7u
aZgrVSS0434DGPU8jSRvRrQATMEczYzh+lgM31zWLB5hMzDkfg0aswOd8IeC4ag4urhBqLo+NoKI
Unl8oZCZXzAhtxUwO3zt6ElvUwQy3tdJiW2554Cu6+O/T9/WUztaRIK85Pzq8ymuvdfa/lfFSR9A
Yg8172X3lS6k9mCeE1V1px76mGBqhtjG1dlcGR8I3T0AInvnPl0eE/KZsrhMBNsPJkGpBbhmNjPq
EESmlHEUyzlVTBC9Zd2LrVug4cW0DXscYTzOf2dmBQ9dBQQOYdZmfIA3+DEnoMxawFza7w39rLDd
Fdmyz9UNDabXTYPALM7aSguN5AB9o2imInECrP2dQVcE2gDBrDNMJ+N7yu7bH7TfzcRN5oFgPJYT
w1CmINdhwsXjZpIsF+giBzrQ7VX9/pbB9fw48VNyT5gfWwfHCalwOFBVPMnInCVvg2uyQp4KC+O/
bZ0tNCHymp2wtpWIry2LbeQEs++jNPhJg53ZLnXqv4hTWuUZIKjl8Jl4XjAILL+xiG7oNt7NozVV
4yyLjeMBfIPD+FjXIg/XF3+qEwSnDt2tS2iHAdZm05Y19ZLXQZsa0fbvzJEcFVoAwhRaP3y+mMWw
YSFc3ldvKIY4pAe1pFofoc30B48MtR0T06wQ44pVYe6d0RFFo5TEa7uPHidkWAoZHGjSmHJKyomG
zODAm8HcWy7YUyh/heflUrC7sldGd6r0BuBncSZy2OG7PgK50Hgr547ONdFbjuOMu4PC0TncSYD6
77szYKh8C0jrKJljbYAN1+a/5BJR418diTdJI4IoWK4FK9U10d6jbzgrxYo+EABgh/Mf7DEbDNu4
D29ngXMnkomUWrTRpX29RPw3Diya1KLY7P3eJAxx5ab+tE1MerKJz5rjEza1/b0iOtzxjoV4IcNH
yj5CL0Q5R16mA07tV4CnV6hKQV6H6fZU/oXhk5gvGIszSCBmP1+WpE+98q3uarF3uD+yBm5vklSU
o0O1TZA2kNVxIBESYnm5O8RnwQQ49+PHk6gDmMvqZfdLWsCbd96JNxtU5F3w1TD70VO1eh22LV5y
jQm4r8lvniLj9ILobXBWJWnEWNYqeVVDzoPbH7McPQY/VUB6hqZ2qu7eNaNXwagYOkA1duBsMeL9
uaeUTo4rkZAofu3y2R3jJJ8LV0LC9VPHfp/Xc8z9Vb0GHfhGq7VOUA3FtcUBSwjnSmkdiWReYm5b
UGOywVmA18e/Vrm1FkigB3a85R+zBBktCSrkEpEcFNRk/SjSvt7pD//9OgT9PelvtfspYzyINBf2
RjRBMgarrI6jiMtnKOpM3xtQ+4HRT4F3kiBimTaSuRhnZtFNQXs4KtTZT7KGB+OrOO1zpMdQc+7H
Bv3g01VYi1C7apQkboWJGFNsIzdgUjfSJxfucLKGBNvGX3HcgKGuDgyIRJgHf5qj0RI6g5kdjYE+
77Ge7moVQpyH6UldU7VjwzsABDu3tFAzL7qGQkjhVyyfDTPj5Yxp1mHbunq8O8wcQtrKu1VeWaeG
QaT/IHJixd0+ELZGzZsNFmW41eu+FMdEyI5uL3JxTU8wseXaNplZq4GTBD35rGpDtsnMYzj/mGRm
1PqGzHtf7ZRubRBcgbEZv0pDslQySR1YsgeAxrQ2VbyOGkGRVscR+pfWfvN7YewhbTzPXgJqkky6
XwiuGkloNdCzD5PGMRfat/4HqJqC2cgkrW8aoADsMlNajDlPvK2qMmAqYiaNPxhZJGnueMCUahfv
/2u7PAvNM+ZRWdsgC+cP9XJw2iDp1DN45izCNjqopnrBE9hdv/VfqdsvLhZPtbKE3wqxcRmuFOah
eejyJrAY6mWXAIcT+0GkXL0PDPVsPmBCB0ST9nDmUCLDiHxAtqFvSDN3Ftzai5+VoliujKa72gr4
mPLRzdgMf2u/GEbrzYbuHZXjLBCW2O7TLnrceKC7A+AsJf21e4jXfbP+zTI8oBgsy8oV3QeyQJ8l
ilMTPfxvFn1MFfpVlvqoBbTOBdOqYMSC3mYFYJLK0DVGLuHTdyH+LTQWI6U/j9r7BZHfSUY/5H0r
oP7sIygrcpJ0Gzq8B2MXwhAy1eTw8lYpxWjGOTk16hQxLIXUhk2yLetAeyVhFeLnYWgsnFD/xRjN
SfY9IW0N6vg2TsDys8SmHs+OVtyyTGx7eNACDQp7uO+NWS0OVfyy1qvKdnxcfdy6vHA7nVNO9h9d
sahsbF6pa6RYBN6xFq2Vl4Sz1i3LAFgVYd2mba4aCdOdfbOJ8OTdaMukygPEvt4a9s8NGGjasXRf
EHoDi4XyIZYUEWr9PYOPewKCHlKgH7BLF1zjdpuK+AXBoXROLTiEOuAZTV+Kg+5Hv7eEGPlHq94Q
gg9lHrP33GE/MhqXuGctVeqjD4Mq7ZtzvOsRJLs7HGPolloegGhTRbjL4orMTtPX57+1wiM/TINh
m2oIH9+R6MkLwQuQPBPCf3DBlHD8vQoLXSfSdEJqVvFWrFr+jTnUz0u842QcNJJksbZuSMZ156GW
lW8WaH7y7Ug+xAgfS50BfZf6o+Pd6nypG8iTFFhqRpN2SAj3CCg7GQrLZ+vliDYsrRN2gXXp3U2D
k6oZq1gy2DuKyLb6HUCqQgWnqNzQplFAgCKBG3G0aW9G7SGH2DptOtLrcX2/kE8ukWKljX5Aj5IY
o8xNYUBU0lI6N9BngSLdyLq27b3dIrBcql9S5U5JLYq9ORWRadf82BVTz1BNVOzmu8FJo4gogYUJ
5zhAbZGwFGh6JL5kBjaP/JYGx57uSy7+F9LH4TI8GMcc3FGyCM/ejfGwpT/RSrgEa8CZPVCRZsnO
kitUuJtPWPjk7wdLz20x1BWpxvIft+GDo3vKp/ffuAHeScd/5CCSK6a4Ty+tdoeeGFtrVVelc6Ip
wXh4juaE/ocuaLH5SwecWecLv0qjAsrz4RRZsNMunwNZ8hcb5X8Yxemhcy5r7B0X1FvLGiuGPU7T
bN5Qqus3I/rKjSaxSj7gbUwTOf147KRMZ/Tmy2DGOXF7OLFJejatIQxPBf5kPuSxX3h0fs/xwgvZ
y/OrnIT57ziGsXjXkpf971um5aNWybOVfkzIol9ul62mklDYbzQMEPoI4WTK02jvAyKTV/Rew0wu
Ca8q6vy6DAvpozgFBznCxjp5b7Z6cLbxKdH9hD4d/GAO9qaEM0pOl6EUZBqxp6krXoqz5BOwGdGh
edzn3t/wvO/InF1x4J8Z/+Lj/3PD7DkkWiNUhYAXzoeShedlCW2SfH1MAsRt8L54fb82u7lQ7jOl
U9zrUKdVaJwpJMCxbkH5td9JgtE/h1k6ev8PNthANhHOU1O1Uqo2XqL8LuY5Yv3LI6uDf/3du1fU
eB4eWL8wFOnNYOuArW3DBOvuZzBRdEtEPU05cRgFUA8EXO2E8s/Aw46bsSugPTXwtGTQSz/MxJeA
viByhfvpIPUk0ysjocCWbcfpmBzsRXn+FOOM8jHfiqzplvAEAsWyE8qCY88ePk0Ojx1//gGyPPQg
1r7hwCaEEyJmFC+hczwDMTAnEbSOrssn+cJEIi0vkDeCDIfdTCx09N7FpOHhFQ7RbI0PZ8I4Qeo7
e1Egm2b82q+HGELE9WpHFtp7vQ6zxbHC5wxD42YrqEoLzvjIQAsn87l7IStvbu8s+QNUZcgyaiwM
1UjKXfeGxJ5nJt1W250IaSR/p1/BN5gKCchmon10vXZpZY9Fv+oY3GijXBKRJrkBnQqxZdLynca1
FwTLOxuM/rXpQ+jEsJkUni8K2qEYUj+3frV8hghfu/ZJfzRBZ7sJHyJXbO/P6YnQGPMTB5UsSrhe
mpQACE61jKLYTyFA0sNeKTkX9/PeJZOwf5lcc7bN42i0pWR9tn8feyt9r/q7EvCtIggXwbxJkwu9
QEgtJh3Il1DBYs+lTct+GPKDO4e98IkDNfyfATe0XjkQ/8VEFBSu25AEYhu48tjlsM/Wg2Snp8g7
ZwT61w3q3SxIQNn1gp4TvKPGzzgm7uV1Pdu5DnypCeGDHefK2/YnY7qcLW4//Mvbl8uRDqojIir+
/aJ2sLc7zbP1zQQOvF4dtMxgogQCM1FI+4hDzpaGuNduMNSHhIGdaUs5auev4xfMVrXh2H1Ij72P
Zj4RfuT62cRu5R/rirN2LZm/d6ZfEsfK3Ckyn92sSgfCOxdMfNgvZG31HK94X8f2oxQ8SiRLywiP
g8NlQ5Fp2Czj1L6VwKcgCp57qWa3o0WOadQUaQClhCpv4ozICBX3j93Vb85MGF3w4ypFxOE7b9S+
O4d00U5icCFlH7BU8uvDBYqcG2B03pGzrOoJ54oW6SMrZeSv70YszNF77UKSqtQ+o/zMe+uin1ZD
KDFSvyuuIB/g+rJpDhH94AiJbSmVRTLgFK00HsKa3xk15UlGRmB+440lcfM2S73JjV5K0+wQT6rF
B0lGX3Wn4bsdOdOxu+y9BZ02q3N+Vle1Mk7CYgHqOB9URXwaVJUB2iqwe0bAi+wQau2Yw9NhhJGb
f0PAIJrSy5LhjAQPTIkBqmL4CysmX6P0UsExNo67Y0EkG35eyU8kTWsAbMVO2hM3wm4uOcjKfllb
vv9e4zuNTRhlMdi5Lg9kasVjCT+F7K89E4ucMBSc6/wCdTgFKXrqtps4eEG3XNlDzHn/nhhb7ABB
IrsyWZzM9v4El+5Mlhfsyr1Omt6RYnTJwK900YHF/WUFBYjHMblPhfktE/4PxpJ540Paoi40O7g2
3lUmKIwng9JKltQcY0kVpm6guM4ZXK5yH/XGjG5M05Z7KzOyuIXhd8JoBuNfbO6mveE39uOL/yOw
u7Ys5PmCg5/2gxKUzr/o9O9PQcmkmfrNk1qmART9OMAwFwpBjvqbYa1izfJPKtCEIjepJlacsd1V
GM5eY/hkSCodGdQ1bKV6gNhNeKDZ00+ceFk2nXvBkPiP9S4Z+3jl2wLaK0RPnDyCA9cfcYlABOwZ
Z1DWlncqN+pktcccZMx/b0hdY++mLkVuNwlf4uyJBt0id3YDWmt/KTp+DzodVkziKuLrd3PB66id
9zjtmBQsYGZ4P50b/jB01RnTPplfryxMPDIQZqvQ7/F3xeKW1/M8QzAvHYPFlaq93463aQR7coRV
+wJjDV2U0i6qCywbCizR2VO3HJbJUQVvSZUi5JyMG4w0GhrqQl6AR7y4GpyaVmraA4JX6RkfUysg
tozyfhzmhCSRqvdKxAq1a91lvnywNJpvxRFU0Dhyn4XfxkeuBYnUEdCmbIbyHlIzw872rytxsbsm
jOyoKAvlepdDb3xR8Gc8uzaQ2Ktsoa3UirLZY9Us286XO2CGe0z10zEULc0hSB3YLTrrKhCxIH+T
RzEfy3SwLFY5/sZGZCqpC57tMj2b/oCZd3jFAmytIg9/j6FtVw389f5tt/xz0Nq36jieRzwbaneJ
2tCEk9q3SipfMMT4WTgBtcmwG6m3XcNU14THyJONveYHkPMmzIMXTO98TfHKPnx6SVDV6NR1MZga
YnN9BshgH5tO/nPVkoaGSo1csJGtxaj09NtfJo0aZ9PwN3XondVMkdq/vCz4wPHGLInveQMyseJA
U8dRA/AidUP5EB22Ds25GYiI+5WGwbonCPzFKCFQlCg3dOLkxe1nazi9r/zFSeX70TfOznKtwhe4
wI89ny0ouSegu8Ht32naeImsaBnpmNwpqVApUR2Pbr1mI8QOqyMa+6MYMwKtoHgMiMm8BALgS2jo
Ujfws6RJq8OPI+cRXdi04LqeiUcfIrxDxaryOJOGzQiwPn+gcWv3B6IqmMmeQnH00KTCmvzPHgL9
4PMqf8TPUFy6RBsOeNTtBTcLX0sd/gGHUpRQyThhE9POLFmuN1NMMCzoUjBLkUCTzyhGADIbqSHh
Gi6uH3NTOyeL7vdPWTnuBdEQ83VkaFbJ0XzC6cXs9phpn9LPdSxOSNOEP0MmaKk5Cuzs/6JoGXxn
NMyyL/gCIfH4mseqixo4meuTo324ZRUhNOOGvReEj46fBNwxNGrV62H9i3+o67zE/d/2AiV2vr/C
ZfxjLwdN77LspYeBSr033g9AiajasYVdiCeuRITEFDJ69i6Cwz3kTjYFMYDd8z3D17RJo2nI2nb1
GEsr6X0951UrZWsgod9l98w256KOFnU9qWheSqIt1x7UHvoozEwE4MWTwuTARsytwalSjfc/Y8uY
6pgriEhoiRbiEqMQITliSjJrxgE61lMKDpR+/dg3v9UZynEDF7tL8ASc/bBKIorK80T0KIf2iQAL
de8GPMYt0w4KgDyZKSw6O1ErEGHWxmkXGNMkUwcgRaqEgRxTZng1H1195eLd/jOS0/i3JcREGnwf
EpzeAZY5NvnKifQgZq1bh6Y/PLT2OhnwWXfggOJQ1Xh+p7Gbhpini4m3r1/Wiahb50Yg+HN4ba7q
yhWQ4UWgV2+ksTRnfuOlmqfqsLz39act5LOQKFOFjvJZfSWsiCjTbYkPnKHk+rEduA5LyXpMgxdG
gKE34NsMIoz3Tw4swVeT03NRRVj30usU/2h+VYUxRf9ROGbjk0AddlHglPDVIcuYa+H3vQBosAUO
14YIkSjdA/VzbPm5SBgiu3yooAWVA6PM3BHtMHEimtDaxxG/byfk+6Pkc+TBbe43YKmqoxA4lI2A
w5w7lY4ViiArYDpQoVmjJSlgjGFUzJxc4ChqgE5GDVJJ1SWMQQDJM3ZPVstKu5JqtoDyL0crHzUh
qYtNCbZ5ZZaAC2aCZ3RVblLsMDf+yk8SnPGPoUyJ6FooT9rf7hufoFzuA1c20JRluhW071Z9wf/2
tibGylJ7sHdu5BAixXNvtLN31tzZZ65c4Exn39xNV5J7QNAme2/kjEW9h9NxjYRQgK97z3s7LXtc
oTkKDY8Az6D3PP1aQr44Fle214bUDKgorODJwD/YGC3R8bG2Jl5FUwagb40nXp2Vxb2haIMQyTH0
zu23DFWudmpr4/TC4VN6eQTeESmq8jv3eRhL1D9UqchlSg4VG0Q9wE0ggwxqiL/ukUlsp3dLn05C
LH0ghyS5Yzo5ktNbUaAGTm/+4LwQL+mHCv6YnNnuMd2y7RMyCX3WP6daGRpOcqMRf6jNq5AK+F3x
VksX9oWtGAnwrcPblumDAEAFFCAKV/wyJjaq3vIPVwZI+cx8y+7ZS4ioB/vNlHS8Btkj6638jZqM
K4mxr5WO3QI99ZUJUpeY0G//0PP3TE6+KrWt2CpWtkjxujcMAIfM8mdY1ZB3Ge/8qhoSOpBYMdvZ
/Dw+bNUZvXHiacd11lFydxXoq4cht5uoir35u4u8K0zb774LGMLNq04OR8bLwfr/dfO6nDNgy5sC
vRwnw53mpO4lnOs5GMk15j+C49KwAf8kY0h5xshV+8Qz2N2U9VVP03+ePO9Z0wjR7v4TM6/2I5jL
WE5zK1nKXsf9Eg9DGnunIORfCeyGlN6lhSol2/6TCLD/hDhekDbVFPNcImeNZCkATtUQUuTfXIOs
IW4dDV2Kw1lTacmWUzhkpR5fVCeYb1nxNNJcIHf6Xg4fYeRNQHGkS0RBzW0iHkLQRzyHPwGUDmPk
mFUofCYaS+QVCLILnEjobDeBKKIiBqqlsXDAwWTLuVGCD6IPcsQi8NwVne0hOxGy4KqNIqbcDYP8
TQx8OhL/0heCC++SYvW6thmb/EirdaiF9e1wMFydKJ2It1cQ69hbc+wFBtZyQ+mGykklZIqYbhPW
kLemqLLkQwPlIEqQYzGPTNczl2uGcLjWFi5c9J61IAi2oXDQgzsHllExUo2yrOsNQ2n7QjFdO+bK
IdzzBVKqMKK1i9WLKSKxEVqBUp5cmbyE4xUFKGesjLOmVGRQBMv0aeC2MwAoVHqhIlnHk40wF2Qn
rTw7MZdb4oQmU+2f4GhpQgKUefQLg1k2fr7rEyYMFhbL+8PhqRz0sX8+uS5AT4oX0TRtnjiTOfou
PLTpVq6ttx/L/B98eOCuwn2oO/z+3iQ1PzRUOVWDUoBCdGrYQO/BRvtPBwkD/5GI0t7sA7jzY/lB
jomXjiy0IVIuVFrJHf8ABHxH/JqvYJHmao5+BxMcwcFX4TlFwmOoswVqqjmQXTm2vNquqh6cpzbm
lUW+2N+XyNYos6ssTKwnq3jAL0C+xsEc3HAa9zmW6R6b2Ea+ccFEK9rXcta5MaszmtqcF983Gzz5
sGDuGy5/q+RDiFb4PChtl5FqbYLO7751aDS+Dai8TTUnBp7TeJARgcE4uJkb3mV7INWQmbAj8m8n
iOwe6yNXTtPJHk7RoraazAyEmvYzYduXpCtRIZab92BPA+xj+RNYLzYnhE/hu7/jokq7jst2d38L
4bBaiO7oWChCPA4xHW2vu4bV3HB6u96dfPQQLLu0kF6ee1Tew4wy/8cGVSwIvEGWa3c0FgTLoT7w
aqhB4A5NA0JeFBm0d/urOYffzXkR6EXV3ecu0XglICh4PgcJhdVHJoE/MWLORZmgbWyVzCRoj5H2
ncj8Pm4jfC2iQbj8sXiLm/sKREFfs8Y9m4RM0/RHmGWcS0zhJuaAJK2x9CQsTsutrFYyY7QQ6irP
Xz1BmSZE/jhI5UA37dOma5hbRfcX2oB1Q6l8YM6QNq7UIZ374zdLI370xCkVzbPU7o6YkzYxZb9k
OLw5F7uzLbnruBmMI0C/94NG+nN53Qmx5hRXsNy5NNmU6D3TomjRtnXeSHJ1pcT1UjltxVZpXgla
TqhFhnhSbQiiAlMyFH/ao1bceISzwamomhjll+ueZrZnpxSPmwB/5bGKoSe5KGRRotmYXZOKv1gM
zGHlDB8UdsTuMc6B24ioh+sWHpq/6smofnBel4k53/peBpYIZ8PZw9PBPt4PP3tEyKViN2ajcWBc
nJIbillUoBYtOtWiUFBPwwHfnkNs/1m3czrKbOsn2Umvkfs7yeCw55dByaIY28yICzGzLI8jjw3e
lAAKTc7j3kJeogiGJxdRPEysdHnXR9DGOEhEK3vq6B4yEWxOQWsjhiSP5JbzvM4r2EGLT1EK2FU6
sTMuKQkZ2YV+sUgunBMQw5QxlywFDt8gXfWG83OmfewiuLu9uoOaKNSPVqgzlGgJGq68ZL0tVTGZ
bUltlCpoQyzmalVy0AUmq3AzKS3DisnkISj9j0cHFjd/l7w7AXCopBWyfYmbnt7xhfyInFc8YSv+
wdmAmmxLqyhpCGp2owenky2ofLowVCg0QruqCvSXQWuY+qJvO/4ViTcxyCJWVQdGGWW/sGQDtDOt
veBua8wVhxKVBvQJGUxLh1XHQmfr+b6M29mZaSUz0rgeeMdG5SWJILp5BQfn+xPKnklaFnhHs+L6
RHZVLjQ+ggF8teF2K0MD3ENMuiA3L2MR+1sB/jAqBShqQijapOAx7KWv3gw8sDUt9QkwZCZMmZSx
WXK8J7kfhHB9yVIsNzRTovG6bcwfAISH+FWEuywB8N0EU+X2fvjKLX6W572gtdTpAD+iAH+n9reS
GQtlLZqnPPHamx/Y+YZk1YNf2buGikHcy9TCPO8k/Ac9Ahl+RDJfw72HXLsMKR/xLOWajKPjOmQz
sLWVk/0xN5O/pGgApsQp7ubDHsy7qdZ0O8H7Q4iFYiUqzcWivxD+xWyorSP90PH1Kr9d4y1mJmZu
OVB5i5Fzruh0QUszGV5Nl7kSX4rxMlUtlV40NUBbS1csLw7f+N4iAOc3ynCWBfSXl3QxgVUeDQQ+
YMbA+uu/DQxUYHt+thDxLAp4DRweggzesZnbfP/4WwGUKFO6xNbQq/UXC5/Yzc7iuyPR+Jbq7eEA
ZYx5h1c05ZuB9Fpz8Q3y/yCEX+4Is0m9Y6ppdWEIs3kFTHqAP+rvd/JhXyJFbqh6OzD4BBNA0UqY
e7iiGxGtV23Q2S9g+Mx7VvYO8zQ/TOYDSvIbxq6d7Bz558pl4ZC083gi40UWbGa17+Dp4UCdqIME
bPHSIIYrIcE4hP5uIHWnKhYbBtcaG1GBvCwTJUNUntI6dXcDUrYKP5gsk0wPwQprs9iH/PT7OXtr
KxeW+3CTbgJ4XLjsZEK6H7uCB78BzobHWLAv8rovkzL4oe/1VFl8n97jXMu03p+q6uOrRkP5GzOV
xJ5/81kR/H9mMcQ6yhqRE+YgvYJRBlNG3NPaozxCzWKbNAX7VE/MJ82mQwnDKWx5h12iZrpXhqxA
uBb9FoHEV50QAnhtl2OqdQpmR4vWflZsU2uEznLdPVucAGb8XglKUEqfL1rnolaFoLKfoTpSPOWH
lt3jRRfstSM0/b8LIZYxMuiTQo8+p+RJr4pT15lYI/bV8ubLqHvLn1hw/mZVe1wLgZYauY5jmtiC
3hX5Cg5ImbqQLMyrXhTcADMvZRopSFIoCUbVJsWKQELacfJUU5Kbr2y5UvuOKDAPihhdMqtvwGX5
GLWOB0UOxQdW9pp8BWSjsPRU6usJZABNhTTHuCkHyEDgRYo89BL/usIzicKKEwRypjXJ+6ZC5gdO
6ztMgPFyDrnJdn6ATUIXTNTQG8TjHQLtjSMjJo8hWWlSy1P/xmQh3TCM7cLuI3D157Po6joRta0l
1fp0yK7l+kERCdm8vR2WiiKGQt86O8otAyN1JRBzipmLJcF7RLTO3IjCm0vH5LFUTfJok1uisNLu
A7hebCnPMW48rqCZzwcUS8btO+NqXZwRxRW6uTnOTqNl6m/mzAWXNzG13lf76PTyP+zoXziQBVHb
UwsMNziojhI1h+Bu0yFf/qeUkufGpJ+gyAFSxQsfsIfO/LsHZq4BzB2gVM78EEwG7iWh5dAplgND
aBD6k7nhZ3mB0nly1CFq83ml+smiw9mNO1C+lTah/KoTkSR8sbVYaLaDtZRRoyiaPeKo5BDiQUAn
WkZ+pHPJrryXv3dLGQMpoBCdrLICjaM8cLZfmVHzYAKgV9wgy7wRKTSWnts9LX44oM5UcpmRTLCj
oUj2XTajcsJqYvYkMZnYGwOu13cEFJddAP4s4RrvrTJ5iDBHurxUj74EhqOaxJ53/QFokg6pnWPz
tn46F6bV8qFQQM6qIfEwyKMsghGHfR6mgWMMzqb1v7piT5qqdxrAyQH3szpyEEQhfvi5/l/vfhSi
sGll2S4gbcuKJWiUDD9QK7/E2blhPoxqJT5a6KgPbjIxZ6BdXtNjWXZiWZMrY1ablwTehoA2pCgp
HnfozPS/AAFezHxSyZ+62p6dRME9kPBpJaFjUTcaJN07/jvpDyvGD4PpqsCyKTuMvLebStxyjaPe
RwhHFHVTjws6ZNpmCtils/YT7gaZaAnxG7J9dKd6qlxTztf2o35Ac5K1CV0AREiYRBov9jOi0aQZ
Qiy1OXDmDWoT99OBuac6Q7YV6IDgPzmPw0GGhW6wdOBQgLlc1sHOK0MJIRdyB2PK0PmjZ0p+Cq9l
faEm6bsuXF3T4CUJqkXbpY2usCdp3F38LHEe36DJt//UBFyTRoAvRVLbjLSajU7eU8vMbfRVYB+v
Nr08c+DFq4U3oKy7+LTC/S7gUGoi7oXUZJXHhgXKsiOKSSoE28TaE4zulObvrU5VDalMIr8Mjj2e
9r9/fBXI966ZhDIACZSONNg7wZXigXE2td+JRLxepXmz+5dgKhLV6H6LOhkEVHHmtOv/wwJcYClg
9XHntclRVG0fm2BXxSWH1cNhl0ZHw26dDoRer4y9mOoPSk0G07GzZSVGRNFs+IpbVJFBB/8tG/HX
ARSqvndWe73/RfeHRT1BSt/DMLqu17MAxWe5n2A6oRl1Bg4Z1c5tcvqUHOZS/BTK0avf+qsYACCF
4XSQEaHqKJNARBqxNgJ1hVsKkgOXOAcangzdzIVtsfNdYyNowaVFhXL1IlFoe/bfDyd6AnjEZOWe
E9oaB33as0upJJirgESkVXAeU5q5zCWOZ9Q1nFmPZEivhk0M0F2yz1GfPwBtS/uT2Iaiq5Q8ScZ+
aYxlhRm8aSvWy2ZO8bUzm0ghCy6WQ2eQb1xz5OYG+9Jz/w7C2xNXlrgA0rKeNlfKt6FgkwtTjqUB
X48yIv3UNTjhWH7KeOPTBRbW/e9dOeDlLjpgAhPh3BDFaEkmbqWZkBlGtH8t02K9VpfkGNsp9Gv9
MhNiQ/Kpz5BYGabWoCgjqFB1gSgnjuKo/i/yfKeftShV220tFPUGitbzaLtYPimK85ctOS+j9gAR
nAvAiZAAX9ZR99iRQbbco3gqAokK7jZqHF+yPx0l04NJzuqSyPyWsL96/R5Jaz0r+5+CfQt1fTni
4DeurFfYwu4ZdBU/+thbQyHGJFfCj5rBh8GJ2ZqjIflfUst9XlTPfwWZAD2gCPwAMkLuSC/ytUHI
yLepwNwD81c4UL/chNDx60aA6CqhqxKgqNWic/gQgM9cunxJC6HiVZo2YgS5n3s0rMprUHRiNx53
44Ih49lFubIaLdMpCBvcQzCCVO2ZrYzYFLUODqAs+RPGGNmJm5UkG0Fzyaul4+Ijlkz2CCKZepZv
Q9/k11rxxqyz9XFTpQ9IKOEEz4EypOUn7dv4Adjdf6qdN1+FV3zmamI4wHzwlkqYVrnVfHUwHQ1P
Otv1yUiRvbdFijbBquuW6Arggbj7Tz577rSL9k+2oeU08kZJxooDVdM6MhjxtVoop4hWvc+rJgu/
QADUOm8+sbFHjTrfEoKnWA2KAtO3exP5mxRayjrdCGFPpMIZOQve3BOwGAqtw7vMqdt53TsjTv+9
5Ebe2qwx/eLO98jg9uhNEzd5l2o2CY8TLb/Iw67hYmsQoRYQgkY1KVjnyupoIMsWZ49Xo/rn7DvG
zc41I7LpAxVJPqrpI3WVKjVxf12mJvWbdfUwDqTmAFA1fxRGW3EcXrFtlExKNq7Ez2vDI4dFU06T
lBp0mDooPFR6wQx6LRnRUZydi9wciYxwCVYOTFvRG2EBjHqaEY9HwIO4UI8JOv0N/dKw2QRafCc+
wJqJ2uieH1YVnZVY5L3ws6bSIYomc9OsmKdLrj9MEF1IGXBpEjalUZozMWyDcEVSeN6aKcd76nvT
gMXPxDbrD44hNODdKRiVoMGw/Zx7ChrWsfhgdMAdFqQsx/sDdzAFFIlhFNZnqNjosd3mKO9HFn6h
E92g6zdhTKG7B1A0BRnW3D13mICZogazMZldqKKjnneQDanV4sc2klQFtrEtJk4QmQr0v7eTjkwQ
/d6WAOJkGafLFZpuYaVzGMnSwh0EkCnb5ObFDZT84YURZyAIFz7PqELYgiyEd6OWWND5QNc3b65t
tGS82G+QYJYGmpot2APDse/u19K5Adl1c0ArSB0CI9nYk7FNcFDMfYntapGW9gf/H8/6coAQSMfD
+aMMnCkyxxvwFtusNjxjITL4xWfymdz+8oErfM/QPFx+6vZ2wAmxKwMQRZRQYve7IBgk1jH4U0Hz
eayFWt3KSG73aAi1c/tgczqjXM4hZWun4XMiFs2UH5NsdRILRx6DgQ+6mQA5ja3uoniKyEphICrw
0zrz55MmmOWwDGLhIYmH/EjzbUC9TfPUiHGdfKrWaSmLlE+AmJm/eFIJXoHG/kf++BpVKvH7q0Oh
3WSRFbTv4UZmv9HpFeB9qNo6kWUGfFN3D4qOB93CqP6EspetLMr+mDRECwTJZqkEvQc3oiYdj1OT
6BhCTRkccymZbLYbr0YIuJR6lEQUBlZpERyhdiMWuw79MVCCizmtgM8ZcLmKjVnL7F5Z548NOPnn
yNd9YG+5QUdhmVbfSNnYe50R5ZV6qGVqrfMRI5DkEtEYBXjSAVAViXtV+toSR1/eDOOHgTcB2lxU
GpexJP6tt/24K7k/xmAsq6nOg0ciWEHnGEaVWK5sEPMS2H3GFtzS2WVCY/sSI+YVaXvdhbGN22LS
P1lDnlCQUPBDGaAs5ipAHsEMuBTn2VQFFKsmbTzkUv2QnaxtTk4AGWoWr4G0zjw7LcYZfxZ80wy+
oyHwFCTx1KvsapFss0L/zphNcLAWTMzr+nhjSdBSvBysowksnsrlP4DNK1QWlLFLxfxNxFrcaIE4
9lPD4Ls+Y4S1F6u40wM5ACY3X8EiWlNi6vi5+X1Z+p/Z/3Hro5NxwKlOwS10OrA22UmNUwQYQVxQ
klhBNGYHU5Og4OzuJAAv3kNZiX2V0n8EfSttJuuva27PjsabZiq8d2mINeNg9lsajau6K7mjAzhC
IwtLZ+MKZl/woSWOQZqwUvBWN0YIuELJIT8LEw9waEMEOQBHlhfNzP9pwlbXpaAW3r4EkBJ1UzIP
r1udr9J4YH4rpJ6+CqvAIM7/k/93Kez1+tsfBrwk3tTIaIpSWU4IeEqp5aTK1a0mAk4cCHD5ot4x
VjAZrvd7XjAKewt++5LOqC+0qzcL+UlKZY2Rvx8kLOZA07sWaZamWNQKzCBnOTPeW3fob73dcfzc
6IkvkB/7gw98fnW50q0BA3QN0fJUIApRQP44YFFM+ZklOyVG8/n5EKhBFcDJ4rZHNRu5s1QU6cyE
lApEnM8jhxYLW1Ui1zXxKI8/jAP++mZRHx8qTiK+rF+OySdHHF/tW2PS84LnbSIbBi6yWwP3Jkfm
tKjJV/GqAzuhHbyLaJXnZKb/LZwwzZ+lVmX+eL/JhjtFB/JvHfNDj9VIq22OSj9t/P5UiYYoTbC3
+kauaxVM+Ys8Pe5EPLIbgaEZuyj9v+JZdRvxi0Jkk7AORdnwY4I/vBZK2lQb8LpfAJzQxMUgn7q+
eSPoCcHd2/vD7Q36ljHHR2g+3Bb71pCRBr1eR++1H3G/HUKt/h7ki6/+Espg722ofWcsmPlrlyQ6
oE057DeNDRSBk6T8S1CJ6TkxXO8rDbidhpFKPAJvkboiFY17xM4G/lOcpdb7j+4hiTt35LTV/FwT
HpaoV9beFcFu7j7NXPYMtwYp+lEO8+pb86DMMVx45VRp4G1fDoxuX+Puf1rZQxyJT4GOu7CYEKa9
SAtvyIWZdKilwqxjGhCOXq7sW3Pk/Pte/k2O1BpOmk3WdU13JJQal0zf+f/Pup/QMUV/7jAk3E60
RSyVSPD6fG5kZ0/SqxRZBnul793aBF9027qOYDadHTrk4e0UT/GS8GCoHLN3Ii8Fe6RgrAOQ+wBj
+E2LcCo4uPeXowaDBxvjgOfe0wyTI6RDNqWp2cCH2SESMBgBkXHRFhF6PVUGU8YutqgJzR58jG2V
SYR15NFdKeBHNKzcSiQqRaXv/j2HZpW6XdCMxK7f8jTdh3A/v+mBC3RjVwvaqBm1rFcgLc8Y8Ack
sGAXNcrR1VetCSjDNWIa2pur6+YzfQnCFB6jXncru1sOYfdkfsSTJ6shJJKwx3ABE3PtEDpIfTAh
NkIIlVIV0/69B80cWx4Cnf6Fo3xEBadm8lQWy5G+fEW9QjbUgaoqTwjiGDiRhragxwxvJyEIQn/N
JYUfxspHush++J/b/k4QnjQfsJyLb+LkR5iHLnUHEsWT93LzwjYEmMya2+PlzbDmhMBSw4quyEOK
hDQ6vpEdOOlDUYOriIBLmCciH1hp20Isjjc8zs9cMmrZumcxqHHn01nlXZEHYUBKjqcXT+50+wj3
6x19Torng8XxKQuRlnYymD9oR+yLYlECcXZV08px3cRwnHXHOGwre1rC1s55ZCYUNHvd1KsSXQ4Q
U+duGAnMECM9/I7wy2Kg29PebboJ8ZrkKpgRt0FTzcHbWLcAi5S/9N6cfKYfY/JlYvMaoMjyH6gY
/vk8RuzLn+cMnUnCUFk57JiLORiBTzTwZceAS3v6xoice0KLnsdHFbQsIDjls0f2I0c7142cnuEi
PpJtAL7jq9pFMSVR5MEA9rqohs1G6m7T7847rN/FNxUsKPHalEZLjQvZNKBncgDdr9+uG2ENNn45
RcHI3hx3d3Ysk5R0mjdrjffTV7ibSczcyXOtvR2r1+rhfDhE3sl9OMbIRU9aig9X+ceEMeG62fJ9
4p4xopgrHZzh4aFyvdj5LbW62lqyTu7LqniqoSct3nYkowc41QLsGTdMWq7w8aKv9ckGtV3xYnO1
B+fYLZWVPWYPgSppZpUTWuTqI0RJyu4AoaXVrp9IyIjtZiztkyL64bNivpKXsqBqfPobASJFbb0n
xSVqJRM2r4K2oeU09uF1+1cgrh3eaSAwKrMGNB+SSrBz1fzEsTX/+UojXDgEVMvQproWVBr0gbqH
8P3i4RywLQiDEuXZhi0Gt9leDiDOEVoS8FKkJgg3AxBMdsJ9K+NvbUSSO6fmqq8sQtsjgsnvhIL/
KcK6YVFfG51TggdXp05X1do1CkfxkYlTze+B6bFTC7IJ3SQJR7ZZbf1/gyEgE08ZNC1VerlOL5Da
VKJuqknU81N5McuaHC5IQ1dw8yErvyBaqXhqIPRcLOwybr4WHuZl44UNQ0BsVUbLEckLLA8Pcc35
MVBGuTsK/ZJI/AK0S954XA7XMToczzI4BFY3knf5X66irZb3dKgIyYtrnFrgPNHGN8o5v04pmthl
GXowPgRPC+rWCDG3AJxCO7WY2oigC2PRmv8fWtp9FkioDNZR6cUDWeZt1UBUfrRsfukU9Q4E6hyJ
j8ojLLdTfYzzMsptor9QnWUBC8XlxNv2GZzbtlEt0lrUpYbuGROYW0zJfXztsetkQcM7N3SsXt8x
bE3+y/zKg0J8EXUqNQyL+P80s/WpcVnLjJ/k2L5lfW3wES3nqcpWi4rnP9TXaPTe99UpFGflgGLv
vd1J46opym/QHOb/g4SDaJMAR3PK6NUszRAmQJZexBJOeu/EAwqWqmGakbhBKK7XbPFLRNeBEqyl
hM3GFG7elBCgQK8VXfnn1ytlAu7kIr3p0hZtqd+clRI5QLjPwhY9sD8i+dgpWAVG8Mbu71tZA7TY
A3KQXfqbDn6BncW2JtZ3prbfHL00oDIFPD1buNAft+oVmHMm7aAa5lhpAnxSsqaCMQRvXTa/wR7L
JrGhtr802Mr2/YZYPK1jZJY0LDM/tK67/d0jdn6t6fL8C17b/G+sQsDsR53XBM5qX6eBVndBniDD
d8jLklaoNstzb/3+vjYmF7QNN7OpdoOZ2UxbQM9WU6LsZpFiMUuSYfNvIPRlwtOq5JzNbyZbaFds
Pp1sGIVXaYyja6yZKulCsfNpbLodnsmZ7Sj03niVuBHm8RWsgGFYbBu8jp8uvLGY37uQIJ2Bpzv/
s6DTdFSwNHO0TeD9ooFgSrE3YC+KZFVklslFJkJh+nBTrQ5w5spvmJB6IylzpA6u6/cucrl68VOh
OAxGgMxGWr+vjOcKorKL/r+Vxrcn1JGKUXD7DaZ2SPRWfxgrp38HhObQP6MSQ8YcJmQy+9GT6FE3
OyENfkUJpeIEb0h28eXiGfK4v3xLBoNE9aNo73MyHqVNiWAeaJAOFiKEuqAbl/pGkyy/XR33m8QD
DLdZqlq0e4qjR/4Oqcc65n7URC7s3+ASW1bdsR9U5nQZmBwKnYen0xDxMgfpm8cMnTZiYXO07aXF
VXgphfW4h81XSxdmPNRNnCyY5W/zQ8p/oYCMnMloH+Ku3CrFm20pfN7VKFjv58DiUqZimebP1Tky
MfcAxamIKIGAcvFp0g8l0M7hodqLpUg+zYufmTyFe+5EiltPY6MCu5plVI21Sepejt+hn30QiW+E
XOj+wP4FH20ENbWX3yrYoWaWQWxtjeIeac51Kmnmy9pTS5/BHDUsadz53T8CQvFqvgdo7Vn/8eeb
/YyZkEPK3f7ycPhHhkvnE3h7qcyogni/KwWC6llY5WKWMAbTaEsTqXnD3iT0XuuaGRr+IC7PA3x8
IfZW7z9wN5LykW+/mj9XCekPtM4jYnpXAnYp0baA/C56sGulBmaLaT2XvcwMxMGl4trBNxdxA58a
PrfMoQQMSoXzWCvqVbSaoZeqXtO7xbExqLbj7AUiS2oG+GmW8APf5RvilfEVUBGkrVDVM8/WjErL
nE1d1aNX6ZdAzEPSvy4cwd1uq+IUeESz6djAq/qEml6A9DDFDKFm4oEZ4CJa30p+MaYbCBikC0jb
S6UBKQq1toAPwpoZOPEpYDw96FqYoZqQu7M9KpIwbB9US1Y5aE+frgOO2V4JkXIxubXW3mKUDWJl
70pD/54ET8SNniyLdqseWaDr7WjTOLyb3zTecvPYPIm4iH1IFj6IFSKoCYKx5BhNl2Or0qiy4Ibw
acmIu64eHo8R0HkcC8jFsnikvoks+d1KI7Mfbbo3VXebGPQkJ9w3qOh38OKO0xFnzOju3XEAnRxH
48zslQE3BEZLH4CNlN/l8w3Tk408z14xF+m/l7WUJLptGl7og4MCpfY/Nr5NE70oXvtLjsQhjrFj
BNTxyVdZPnSZMPQtqGDiYvCAUsAkW2hpOLm1JEg1CCwA+X5SuZgkbIsZYFaapYGOG46OSfZQMENG
/03HymekzJLiQtcQ/XoHYtQUur+KYdwPGPUE10rnQq7Gwhren8VG+hZ+DHsLByeOJtnL4SRwlqQe
Rn62IxDbi1wsesqwHD2aOxS9Xc05vo86VsE/h/NJwqcBKEJsYQdy4+cYnjwuD9EFJqBBRvvzSDgO
dMletNkz3WtEVyq3MbzGciVB7xnjtEh3XaLdTT8JJhGbO5qQ+AQR1mtN93cuwN0mIUeI8KxGN5oE
mLdjx4PkL0pPSr3Iol5xN7MiNoqfMFQ3LSPG2zw2NZ0EHuwGShK6vfqq7lnSTzvj4g4YctuMJX3q
qFDHyu8jwZhZ7RW9BdbPmX1ZQ0KVbE/DDN2ANP1Hd5qBxeOAg/r5kNjwHkWAOvEpi9OFq9zqFyVw
3AVSv37zojkSNPoVnj9EDfmYMsRwAXuzWq7Gzg9TJjk+eTxQG/80CHwsrVk3iOiwe8ogoD6hOxl1
bx+S17KAfRXS0mO8qESMcpuiE5KMyXf40DD1LynksMFjNBZbys6odWCMXxabhmIXCppXTmVEReXq
yjr25CS6PInc+G013aNkOwYbKLZarg8dewjxHGwURrN759bHQRfK0Dbcc8aXQzCHp/k0TY8rtp7x
dQYiTemK7qpJL9hvozZUpFd/4NDkZkZ/Y2Nwp8+TZ9vj0x11Hh/I+O8fxCpLXUwVwb9GS7QvhY9v
Vffu+4pJbM2TImIe97+YXTEbZIcxdm8vDpoGBWrHuMsP66o+yCtCJJkC4j1bsAC9MafSPQhRIMIh
IfNBx5JAoGjyd/Y0bRuhkiXLtQ1OlHQVb0gR49KbU9H+doumpy+VYYnSsSKMgjRDJytzzI2QKV72
pW13RQRKjhNBRlnIy9QHy4KJATnUdl3UQZVYQRkXoWWxTcClZxa24Y2PTii+A43/juTFEnZMmvRc
kXSJdtP9hrv/URoiFGrWg0KKYnKEnccO5Q6LoPRMsArrrNFjddIWwvHQ+vMWN7nj/q7FNk7iwde6
j+vbQLZBh6Er2Tj5dHaRTLtOHTrOrFnnS0Hv56Eh/GRgvXV5bNqGNbh6mtCj4TuaotfWzX7lzKO8
zNBDppOWfgNdrdkTrvyfEHSKz25Q3myTG4yb86wNCJZetuHEWej/c7ja4K6VdFcz97U7DZ2P1sQf
SnNU7UdQbVUSyHYIn7YCy2TaDUAGa52qGCKZd7cnSrOKQ+/dVIzKPBB7x0bMR43JfvtbdJT0pZLl
AfjUkbF/ogyTtrVdysIIr+pPBEsG4ZvCJh0zO6QBISAyHTblDo/pkkfn68iZ4faWVaIJrstax4D8
xhhbx12iiGzhAJx498gwD7bcMUt8yCP6i8ouS4LThRiElOpbD9BYThoL7aZhOwFk1G9zbJKS4nZ/
jAgaoas4N4kFTx1KW3Y3c6vRM9Y+dudL2kBf1Glhe/a7vNbz4O2z+/62L+i0nA5W6CXuH3BDsn7K
quaV3O86e0OMtd22ZCLP3xpT0qrBznxV1hk5AEWC5eSbq3XRCxJLfsJl6GviwJxXBi8QA0DNdT1l
UqfFq8sCdmp8i0/YjCGpnGId/4S2L4Nw8VAMVyNPiuIDm5Eyyz4795+pxIhqHxKXDO0uS6hNO+xW
CgcREkSzHA3fMvpFTB6KYnDhEo3KbkbP3q4CASuyL5KbM2dPoSX9YkQR87zhD7SMNGevi7ZmFD3p
1q1zXO2vm79/jnmpnBOlfUhP8bTkQYRgd6Xc4YW/zAH2bvLUTONpXL2n9UHzsPeo1gWsRaO7Icgf
e9UyW66f1TXUiYC9+L3tUG4QTjuv4E1GeTidTBSxW6en5kO9JskR3zwzQUcVIj87GCJMduAr8BzF
5GskcupUo6ffqkSXrHIT8IQpd7TT02selV4wSpQs0MxtCUyBqDg8XaaMIKmfjLBdfnazwfYG+/98
dkBhWVArXbR6G4AsZ1MoBbrhimOF51VTwwUcSvQS8zvrd5JmU2SnvNDXdSfsX5w9S2bZdLq9UdZ9
VZsOMYiHfnhAOYf1Q+BxpUuiTt8S0UKFkq36VfQZ8wNjzF21M8AUt/xtgy7y1eHGlFAqkercFPH8
QrGiE6cNu32kgjPZc8dNauBVU6k08p+MP/lOPWKpB8QHCuh6ktR2BLOfr2rQVwAtdtNCg0oIkmnB
J3yxjBtPvw/Ndp5dHbYgBWS2uzJ7c6dNwoMLI4WAEDnXvi4KkdBcrcuVZJ7Tneg4AhFHdt0AWcZ6
RqkWiiAzlUPuqeWHbEbDr/yzOPeCx9O4UxMnAshux2jeY5+Q9vadvStRFMxM9PYxb8o2IDi0+8bP
QQP0NZTTXI+HO5/dNoLqw4JO2bXy65FycYV4gMRSTl1sWI3H1BjyY8tXbOdlUsh1ve3+fnlZr06I
b8LigQjeRMOUw2QA0wcrfGcB5ICcKJsIbr89RvWnDHzVWnTWBtXxerD4VGymgagS87ZaESL5+A/b
2NNYPvkb2l3HSvw4waLVcDTnRUQnGgKWTuHv7DT5TeCI5p2EkqwUGMNvq6MtU88qq1RPzqW4Tp8e
ZTLIm/paSKCGdvvEYAPhJATYxPk6dxrU66aHQ/KeSe3IoOm49hk0wKqiTGDY79UqE9hB0aNZMnxA
zLkr8NO7AX+T3in4Ytjp3bU6bInn6AtQEyaBJZaRyj9Myj5r+BCZuNOYCwT9uAAI+R4O4CLzmRIc
sofCqDHszrplngi5jFapEGKFko862hwtHryOFSHSBCaCYEUceew3wBFPDDlPRYFN/+S76PPO9Vlt
X0KultjqF+QKrzUIJ/51SuOf7hy8tHeg+hwHBJU6TRsiYehFHQUa3j/tvJsFGit61o/T5pt8CTgU
v/J+IQS+DuHpf3VTyZCi0JHe7pkzSEBeRKR6YSETh9RPfmlxR916WxhO+EfdtydRtb5l8icQGiag
R7v1pwYPEc8I6tdGjTZYB9BNdebdyE1Np1GNo7gG7E73BdP/PSBm2vVORSYXuxwXvGQ0JgUeZB6x
/ViZ6jOQoPzCnPGXnX+WdXXFUe9ixU4duLpEY0lhRv9+xhTB0vVDR4+/MjRK2NSloyrbsEPJERrL
8W8rLFb7BCGoM7aIFPmY4WqJw6UlsQZGrmdyS9xa1QdR2ubX4N+y80JJL0EvEaa9PMfgsNrShKPd
OmweK1ChkNGjqfr1Vs3Uy29uuFWNaeoEpgEbUXylKhKNUfgi2rnarfr2U8E+5kFy49m3feB4eUyN
vbVipF3QYusrUtdAXDbyvSPEIEacQiUDBT2kIJONkUAnyAgW6yenv2mn1CaRXvTtZUoUnR3qNz9/
1ce8THFbbuc2LApH0VnfQudectsuNaEmAYuwbayq0T6juBN1BZwOZYRAu1l4P0RnGY8ff6U2HSLi
if9DbV+e5VUoJfNvzJdgHBrafyUgG9AFAx/9mE3Gl+qN25bFvTE75nGLZgjqY9SbqIjU7sJd9+k9
EDagw6MKm2w2GYCjUWHTCYWQEm3bDug05AHx/fTkQ6tDjJKrjsCabYLW6MPGUHunHwoeFXSlPZz/
7J1GXcyD1gt0AODFfG7Vgs8IF6n7ZGa6L8Bw0fAOcno1z/RByjeb0jxRHTBdbeLKUmpPIBog6siJ
dY/N10c3CE+1LACMfD6D9UDqGyJ+7D+QTMz6lPRskYu3UJxqxJKYm2DvccLhv/vSBN75by4sbBL8
ks3IVr1uUhk1ubSm5vfsN2HQymFfNl/WSKHQgOXA8THob7thtTU9cmgvk0cdLYYplZKZCKU0NqrH
ej0LLc9a51JV5PV2Y/Shu7AKqsapwb/dC8GZX7qGRIp86fVrfN6GfXhw1I4zW14LUBkz1ktnvFZt
TkIyZzmW1LGxGVi9UXUkB/uGhVP44gGsNgRk45nF36oK5s1e71x7MclnXJIn2d+Xz5BbQ2QuAwBJ
c2FPfU7OOhhFsoeMzrPiy3ESNry51uy6i8XujUV51tMCdHLQCFht/OmjH+CSy0ZPdAT4QmcdJK1P
i+opn5Da/oAOM453cLPgghw6LC5d27e2MaoWYbUFH6HgR4tEy52XZIO+ZtCZFNqZPEjeKf8EhBzX
cqD7jZeX8Ru8W77F/quarhqtAVd8RsahPWE6jMuyqHv7c20KvILLRw0Vz1c9Ove6gnDnkF1l9nY0
VXPOg+n/nQQyskoAF0zIeSambLs+QB+exKGEYo+dhiCTI4qEGR+yqHjDjTgppP9O6/QAPFS9uZBT
5GzTvCBiukMWF8sCDBX+r0NEDfiwSyf4sNiyxdy6Bd5LdLRdx7f0GJ+VxRI+joqONN6gSaUNzi59
BoflYHpsRJ6nY+gGIQnk/3+QHCY1Jnr4gskYY7bLKXWGke7DgmwQosiYAUvqnVndexJZXUovxpGL
MUI87CtU+5yv+l6R4eHNSazUAgtb0fjv6twzJffXmnxgmO8Gr7cuBN5FudeHKOnjs4OuHDLKps+a
2IKvqPu2uIdL5WtWp1tgrmCG+pH4ITY8sxW1BMuEuJJnGQkIXkVfUxi5BJfGRXHYM1rdPMHMZALB
2Mzo36PQE2vJJ0M8fZteEW3WK4OKz1jL/WsPz0yRKKGUVDSH2dwOTjfWf6FZJz6XiHsJ7l0ioynj
WbIUy0bVnxooj/VHDoRWdMJ7ukfg/Rnn2m3+ePKrzUX5WSjyOJQyC/6DNjLoQ9spf9znDdlIx/oa
FCeRWlAquSgxDmcnxfUN/VZpffhrbA0c6uEAuv+HuzYwPw2QkMi/1NWl+DYv+ZaNYrJwdP1h3STg
CB7UHhO2eY1kFz5AQrWm7TPxvS2uCqt3YJ0ZJ1zpNHG1Nd020V8/8rX5tpOGUCJ7Fc+v/ESmexDM
JoMFgihRORys8hexlx8JZ9milc3ayevgXSouFVWB5mOm2wIx+BI5ehnHlqx8wMrhg/2BNvSTkCS8
wqEJp1yFtybnfhmd0foB38nAyncoAeJiFmcGHj9PFJESBwgWnSOblfpTJXoQIkKcg2IDrYATsgZa
+Ia66nBXFFAZYnlUj1txAUsGq3bpku+MBf4d3hWrC6u/p0lHD8r8fcrdcL905zWQ1XNlqJFWVwZJ
d0aXyFQiKm30lNwmUeVGqud6mycLl5+o2qEqi3Nc3UaPwGnLpFQ+Fog3LF68MCI5b8hJfhCLaTSj
xbpL1YjppnmliXa3Wifl4wJ3j5sE4Vv1JRxpFWeJq35COnG7+/bVS/USC5o3gT+KI3eowaLVNGlk
HeX+Mmy7zDzNeVoX38w7+fG7y3etjd+3FS58jXte5u4aEsQgmpP/SzG9PqHsWuD73K0pv+yoMWt4
I6PGgvSJV5U9r93pLDKo7P1sHaiCsxjXUgpFX0cWe0JuO/PC1A6Go1Byg5Lq9RSplPM5+lOeIi9Q
TGTWGYBEjfFoX3onzWT5mqv5K0MRa9r8t+0d4uM8WX1qC46i/JV5kLOkYVc5NxURFtmbwGk23iwU
I3A+ynuEqVOcaY1nPR/QzqSa70kHoeYXIaPCMHabl0ZUztNcAvd+AzXlC2C/LX3Ap3sxJbfWDEL/
7RR4QpLN7Pd+Tl/dAFkvLUjMa+G+jVkoQ07oixkYfNu8SdK9yA1m8SAvGFkxSbaDVrGdmAUXm52e
2cSigTK31cAj1riLcmWIrDkuhVNkfIzhSAODM913Crd0UuZVcoHvSEuOrD3LuBZUXL2XjkxeIZZx
lLIaQ8V+xXt3R4GBd+jNdKjU9LwYz0h+g4LSjr3fRtR1Pu5xUQDTwtY/5Yn06WYCOd6yEhni/Uny
sd+8SzCHT9punMWTHP/H8X/MFsYlxaxSDbdkkioa/YrOs5K8qsSWBGAm4dqgR0wBVx8ab4HZqGtN
TkJPAkda1a5CZYTEukkUDX8yLXlp/fhGVGm6QXYQIw48QNfbd1BVNeBzAByOElVWOlUEUDativ96
oaHbUvSFCmacXAGQCmgQkCPOouFbIWya4l95LU1tEhA4e8ydzwtIYHeyB42UheUQIRaSVJQmdquQ
FeIUEnJpLolBAj05bLaiNMCU9ZzTa995lngXYs/ItaExY862XWaHBEVSIXfZZaV6GqdgdC+T0q8d
fcm3uQAwoJvlhbSvhveH4tMWiuXqKIpxsYmXivgtf2+TsxHevIxR8Bqz3oWboNUcyZO/IKdjwdcO
4wda/UlTdzWOe71xCMPPjXgnzU3TM/vSYlHrf2dt8mpMyQljE1Hpnmvd3lPBPmjB8f+uRWIzWApw
Tdiow2XS441xSejnvjUMGYRtPJuWvU8IITFiv1MAuqEUv/Sm0YtVBGaEnwmnP+llOB0D8pP7MI5c
pt5gfpaP/jm2I2gG2TmRrEk1DxRfuA6qUp1pqvyKbUh5SBJn8nrkSFkpK6r7aIcIu6DBEnrGu1Ap
t9OGyT6YVRH2tysu/wE1uiz2rZaeRYvcY9K5teB+Oxvefmxsi6h8UrPmOtNX/FGCcWxEymSN7HSk
oDuDmz5d+EcPONqbwIKjuLxMBQ8ZQ8LpfFu0Tygi3PTN1evxeZ1qfPn9Mplj8ndlk0S1hhACJa8I
npsRIKBfmYRDVyYQXEVk4VzepZsW3rGWl36Ll4cMeBlCAmCqUYlbQKPw8uKG3vOQPf/c2WbS0hmX
h5RVnX3oUwKbzKQzaS7N7Y9ts+tz5vdxRRSbz2qWBsung4+J3seds4IDt4BQwiBbDV1eQ5DBbsM4
BsWUPW9PcOGYWlvgvLmgt+KtWdt/RVjxzfr7km3N4K38IL1AQq16r30bWv3/WB4DDT7Y5BhCb7XS
xLMi3UZgl1WpRMUoXuGqg5pi2T59S0nwppduF88y0vMyXUOGNJ2EDVDawL4y6e2NJ6XspV1fp61c
fWcWSy6Zh74XD68OIdp6MzbToMbB3QjVbVZI0sGhQJ0tCg0xt84tj4sVdJz6oBicUaWJCGjSbJX4
eLh0Zpvr0ak8hiiHkvgnL8VwuqtJFfPl42/RAylhFpPWJxlf5pR8VePbEZXeSPzGiKVFFD3hGdWW
XJV5Eewc88vQURpbUfjY1MRAPcuuxUKQC64ccOc9Z9h1To0ornI8S+Ame0+mjqLRV3M9Vbg9FndJ
hshzOB0HbJMsULTutzN/tne3dAjHcaUmQDm5mc1wD67a73khcPuLVtO2UEiVDl9S1zUUyKK8DLfD
XYp1l4XnwBBdya/TzpWsA656rpxi2aW+RWCM4UMmlLWJBA/nLsX0OFBeI8hfSBl1Arrt/VecB13/
XmLhyZ8pYpBoDTTGXrQ1OKRlB15AlQoxzLJlpARrF3klMXaOX5GSJwLVU7Gt6YkApKjIrCsjUYXa
+rqwPgTn+izH8HprJmzwO47WZMkB7k6eVZmB5qqcjbj4kARzJRELYwEXFFP/CCNj7wcS+4FLzuuy
ea7B2G0w88h4BAz0gI8EeQ6MvmVxELNYeDzNzlXorqRybKNqPoodNAYLd34C7iX6I3HxStD+DXG3
bZbPU8DmT9ks+WYLGs5tMAY2JqD1hsTs6LY+wCFrgOIds0MnzrkeOoDzIIWbEZAvEJMqTNfaAD7o
CZ0aFNL1z38VUYIUfFTTo66RuCHi2DNtibptn2Nd2Buic49X2PoIumkJ2YSTUks6BJaAn7x0BulN
iU9HNs5WXAS06Ke3sFfVBXCDUG01ssY99gaj6i4VGRUOmW1YktrAyNT54e/g/5Z8dwqqJlz0hNNt
LX91uaswa+sOgejRqR0/BPQGGnG4pZSZZ5QK4kxU3kiPYdd1A7GNGSZmEW0DhwHljio8adDzEcOa
5GDVoI92F2txdWhukvIiLcznqpECFEQXQVRgTmSBk7/7KPbmTFYM6jdKuwQE62YiLi5dlpUk07Mj
ejyeW/qjtBUQeWzX7mb5uPFMhUC7Z8Dx82Qmc7+kSibktkvUEJXCC6nUhsNkSBhD5J3SiIBSOvew
D5RRLvsz3kgrWl6UjLOlf2CaViAH8tW8Gix9PRSePvcdM/TyK/NaOhbmjld9ZR2Ymnj6b6WNoyHX
SOHceF7cmSaRGl6rZsWxIhM5PP+m2fd/yWVvFBn5LsuHQQR4mmcR+/kBfKGb65EaBaczttDTmu5B
UbrOBi1Gspuk4LbfSTyyWeGcImoILNvw+doIN+QOcKDqi2I0C1P6S+Oh9wqC+Zk+EnbAqIMDYeJu
2A6y+16KVe1SKf3cEHZ4aGuuUjlWCoTPO2PdBv6CWF+HbGnUjwCi/FPylGLd/fZratkCbFqNKF6x
m5oGZxWmdovErsaPUhX3B8zaRL7jiKDRAVA6rIvgvhotzv+2IU6Qu1Rb67XAfoDop5FwSSYlekt6
cK6b6LNrl9EYJw8evOokPlSCJdvh4b1uXqrX5hF5yC7XErEp1TmK7g/B/Sh/YxJvDBk4qzLd4qjp
IHbjH21UxuEfhLKfSOuvgTbz2WZwicZS1+6/7jBZiCZmKLUrYRetepTXt9CCT9hoMW08XvDSmMZr
VYo5smeoH0f1FCbTX95Vra0F/ItcKUr6jKjP7ACkniuTPlUU6Eoo+/DbOQbImo9cHHAIRNnw9VB3
xC5EAev5CV3JStVcbUrJWm849cS2phYFacSN0IVeUPO8ldh8o3Ju258zV0tFYvIwRzDiBmbOPub5
nsMBwtuGTfvfTohLXfTiJFl2VfXvVoepUF9kKKoZ1hMml3MoZY4Gw4YiFczEKYwpzyMcvnb0KeAe
ByrMT0Y8q8U2yDqecEywQOTrHRNAELbAR8T+067PU+nvAx3YVLaugnFjHYaJTiMifSzszNlEMUqP
fTvmTSHI4DX4vjFRnCXZqSnpR79A3MjQRN948EqKa5r7F3+0dlw3Qf4g02fZZvipMi3E5/ws9YM2
SxxfAITWCvIaEGBOOFcG90QuZ5lJlOseQUrXU3Dg6ZfgkqPeVKtT9vHvVPIjvq5ReBrNxbvzygXV
xAcUg4hgmr11U/JNjyAbTDJ4nBMncUKh+1/EjySsui+BQom/m+VpAGJgQOu8KOfosQg2KT6Y+WSr
9gDc5lsX2D5nJIRU9tEnWyEUt0U1mLK71aSLY6ERdmmXLlFJkc+Hxg9YxMAQJ4qQvuyfzY2bfUUU
8aRP6aHNqWMc8IDLmPwi330e/a6p/lxd0X7oPBFgp8Kdjl4MO/iFezNQiXpx2xTY5hpfzIaDHJtW
xc+ZykajgLCVusapttGukTDL+lgK6vVzwr5i59AFSJT8nehiX+gXcT7l9NJQt+bVzPtriKyT64Au
mB2su3GrPiAQmhJaa6/saNhNCVEfUisxqDBF9WIrUfwVLQgwEa1PDdrLKBIvy4fc8ubAh/hwKqLZ
POK6Dcw+M0z+FdvIIRLWndustKNmic1JgiUcr6dXFsYjH4zsq68pTx6sh5qPOkJVDL+elfzGbUG3
+yuJmcTsiS+NLXIeTPzSUar9sYWU0+AEd0kaTijbYZMS7qVfm8XUQ0yAwfTQeAeesRWGTxCsw9+4
zWLb2YJwr4ZEb8X2M3h1wQYpnA7MBNJeDmLFUuKabVmkB4iFOq2q1XoQKMKlyHnQ/gyxiCBhV+7o
qxCcC7KgD6PH2GMCtMg4lFuelKno34mGo45GxHpdgBHw8iPvpsm+WNEVnKAMJmJ6hFJjLWtr9Iuo
1JbQe48FuPJ6Md6FdO33Ischf3lMZB+HmE1znlsH247EXcY8aMamDijINwJszop/p6kz1Y6LODsH
HzyL9b6tlm39Q9K/Qb4S7ZnciTflLIemBBo1acxGp6nDgS7yMr6q6Gis2c4hlHKBjtdvbEoSBDW4
h6yd60QC7t2EvrDo/S03sMAeg3FoTm69jXpHfPCJ38vaXUDhnvobXxBLkJzc+Nq+2fodI+V5gIdB
DT0yE/HCK/eHk493NxWfEpyQOk7j/M4PIqnwRnh/L64+vt/Ob5PVLwhKr95Fk7jXFLMN7N+F3YqU
GbNTdi0CWq2fqfk/ls0kncZ2uTNGsi+EhWRW7RVYrpIJ4L/mEdq7Rq8x/JpUVXkRLgGU5dt5a0S8
SGEutuyJ2a25Bclt71oq/Ezj9H5qRtXjk/LmoWGXirEpEaAICiUgeQsHi4wuMk9jnBGCL5hglPkv
UWdk9n5POVsB4RG4nJ6ygy3MThr2k/sbOv8fpUiuAO/ZH6B3QiA1uYAY6z/heGqsktP5MJNx4ewl
uT8u4MRfY1sV2a+VqZS6q3kFBdhICciDBemLuIy85WvI6UbQnovepqG/G+sJfxL0vCQrjZ+rj14k
0upIrNZeYO5ryDSt8wgaPQObLGnAWf2z+JaaaLd5566obRga9UZlmHOPfPZ+rchDyJ/oZpx4jWj7
stB3lM2C/7pq8i0K2wEcmp1UU2ZQ+xf7VDZADPu+x8oZmEoct8kfGo2IQX61cMOjGJItpAsSLk6V
9oswA97OVTUPLeFqDCmvH+XMUspq8typ3Dj+5HLWjJ/9oRTSTXOI+gpFHavSAaB4ffq6ipA/2x/f
DKWhv+CIahmT1Mk6NUNRjN6MQi9pNGHyuavC+JrYLaagD7K3sJU6TyGzI3v0L+uCrxRv6k/KkVxe
NsWT0kz7q2qPirgpDDb9OSC9cx5vfp1rQWosxvL+ixaKFxJ0KHU16puE8tywqoSPMBpDBFKaeZz7
BbklVnago1ursaJb1A9Ah3ITQ9UU7eHd7GRi4EchRu2lGPoQxwP7nh/KQIfD4YJ2TINNLqoilZbW
Een/roqs20AGh1pp1jyBMyNoHvOqwjvxmb22sg90uSuVgQYz5YtspE6LBg9JmYGoj81Cr8atE3uh
MWLWG7kvwBex2MteQDg+LhVXbroi9asYF18dZVH/2rKk9IF7xSuskqXvUeTntak73iUFTLiSJucP
KyJeHtt0DD4wi2EyRF+h/kIBBBdnoV07doJwPYBSEqSz65NppLkRb9x1fbXZHcItSFkoxdZTFEsH
/uKC1FtUmy1ipV8+WwCNj9D8dgZu+HI695WBlw3HthUl8y/fZxOQq6nmNUsmwlzcgbBlIVgY2Xgo
2oLtyDFNBtG5vqtn42SfUHtfV8iimcerHhY2xXTNgopMmC3wFEP07jUFrmGJXyV5H92qwFrd8kur
D9Y0nNGcgfOOB+npb4FTqlr4KU2zFFWjICnsAdXsEtPy932aiSJ2BxoI3dwW92X7heySElM47CoO
FPunz3UcVlWWN6czC4pIae/4V01eGgxRE3YEJeRrks9pNhlXPJZjmquOImhHtUonOcmcf7tUmskU
ZRnqFBEM7dTS3DrBgvfd2QjJSCGuFlw8uR4IaTCz5P04YErCem05R6QTiKEoow0BNmbh/jRntqat
bTL2HWfRMWk4U0D9ma7L0mcjQnrmUjVw/CaelTAfM4TdkjtVJ59aIvmxTgBH7/dxY67ECpT50q3G
yLNwJiQZpvQtKa3+5ScOWLOeLB/TOHveiH7uyFG4Evo/8xRCFaC+zS+TOmr2I6BLQYwUNPOOiSZk
17Xyo917hWwipyi+HIxnJbTZy9/HbFEyir2FnaeyOZ3pKp2rQBVcYn8YLNEIci+3rCcxBWAchht3
TJmq7DcS9/OQkzvtF/lc/EVO2rKQeze2FNLwGdr3DrNWIFUT/WfnQecAgHfnJDM0ZpO/k2bcTH+R
r9ZHSo7KGHkXjL0i5JslL9DRiTGgQBgB57i35AUt7GvwY+J41nSlSdUPkbzBYAkuVVLtlxT5ZGC+
rVHJqZvm/sFRujG8YIRkz1wRjGnresrnxjYSvOJvt4rNo2DbKL5rQjbID2+qpwCTYXHNPArm5nH5
NzW06+QKLFASrsQkCiZf7rqsGjHF+Ymzd8A/zKEhVvEbOAGSz/DWWgFD0F6bmJ/ULHbyvKuWaaES
1HSaNbHETTjiztfYMtot+YpXBirBukmPGj8JNZCR7mCl/5pGy0FW1COVXB1QVb3olyDCMb8gZ/Mo
Uq1fx4P/Jsyxon6tqPILNeynjQ7GBtXlRWKTBJDD/2hvUY6YZ9Nw/9FaEKLF/XEhACJjL7maV+3J
XAtvOdUvYsGOR7y5SaVOoWniBsfjCVXm4c5QpOBfz/GUJolVGlISh9rbiJMVrviKraF2enjABHNv
pt/UsSLtA2E/01X8W9EYDcI5sYYvt/tzThLPhvX/9qNG/QwEj2PqsN3Vmpw7+A2E+JFX7GZyPIDZ
TUOcO9Hd/Ak8J663BkrT6mLpKkcm6yEgV1Ur3Okigjlz2b9z51k5I03Q/coH5uDbBNLxdt7t9NPx
Wi+TcOcMPZz191GtpzgO/2hg6rvTEVGh35h2nNeDqC7P4SdYGnAKft502XgED/cXkXPMUSjNKimg
6ET/63DZLyz5vJTK/l9I/LThktUZu9JJNexM6zNdO8aa6LwjS4mptoo0hQTda5PZ7uMVu/0uJvL4
nIAvoXf4Z2j59ibfeHDOcZP14oGt6jZkhlztj218oRrziSv+WowtHphPTG5pagh9FOm7mqANTbQs
xiOptDuc6oPrO1GdU5KDIcd6uKqc9UARlWA6oLANF1tpMnVKCg2W0WvgYHYUBM7XgoDF9Xx174kf
kziizXDhUy7dkRSjA3qTZhYCDdeMGwQJ/A7yQyI1IvPh4jGtZP/f2w1y2omWPrpY+k5gdHTRJDwg
Tw7NwF1R9BBnu0BSxPCB6I/GZ0V5baqdX9ri5PEfBhmtg+OChz6FdlWH9fi5YL6fMxPJ3Pt6W8i+
dC57JvtYvyOE07ElfwtbeCPt7SUbMJgmV5XS+q8ZiUPdtQbwJRWWvJuHWCioyfFP1xrGCtfSazS+
/mB37eovOvIZLugow3rX7vUsoIbXrYXdxANUxA2epqt9sgejBGWCs6Ns5krsnkTqSZC4rHT4kNBi
jinFYhE3Im0cztCybu+ZlLbTAsYNKJyLyXfDdgBzfbYFOFYZv7WFG0bV2LQVMVto4d507b9ulDoj
P27HrkuFGCXd8ISzu4sXPcEloF+C3q9EE+G6GM1ZdzunSzksbVMqsehDDsnT+jbtYznLifWQMgBo
rVsfBkIzoeaGqAcN0Ab0IfoWY6OzmiAwa1ZTIqEd6eX3ZmjUHBc4LmvlRKDhflYPV4knX79EOEMY
Fviy2IzXOm918Qcz6YI7F3gkybjbxHtqLaWLCoEF52CLoeTImNoxMx1p3c9EIxBQpFxmQzWL8JT4
rZQk+bJ3iYwfFJPHSGcQA1sYwWtXcEbmHbaTj/0ji4FrJ3A4kpEHbsk5CL4dIgKJNXeHsg0kg9NV
WYIUdAgKr7E3OtTzpT6sNw195BYbYxv8gNBcHCZFDawKCOhbZgvvA6evK7wYLWCPoh3ZvcNYxfSF
8xHBRR48CzrlN7o2mB4awP0TERzVaeavdw/Cyv38e8t2XPb6NQQ6TivKflWzSvFrm1LfNA2DHrh/
/1UpmC/MjKl15MQJDt7JIh/qkxgiQTbnIzzbWNx7/YTbLkKEGrG5+FjhZc7AxyOpjVKHZEwzUC7S
+6+J+oT1+ufXQNWMdeEaiiZxFPDIhTT1WxMle+yDqn0uknWm5C6OzhrfzWJzEtAz9Rpy741TrrL3
Hjfd30Qxxm/8DjclkvQdEwKU4CPB8cE4on8R/WTkbOSD8uPPROxSF/jLJk5P2R80nhOFTVf/OFZ0
etyCsID2Sb0oCo0y1xwGJIx5NnXj7YoNEhPh9RhEUDg/ri8aRP4XvBplazCQN7qnqANj9e3dGYQI
9hVCuphw718dBXe2XVhAGb0WT3fEfMddNSIRt1VLcHLjzcXp3xOuh9t8m0mYqJBRdGftCskoTS9H
5DFCfchOfGUjVku/t9paPNGm1hwcVuTqtKyf/T+CqBt7MYBdpiQcivVLW7sBSxbjKn+FgS3DBjyK
VfQOjs997Ddud/+aRsVmsrCDU/P/0LXWPHahBkI17PKWb3pdQob1bo3pHphNeUQwHybrWwfqeqFB
hee+TPuWQFId6bjwMlCp6DMJcKcJ0N5O/J3q3zCfGc5UqvDCGEuu+yUquqzvYyAetkvLI9CPvwMx
WfH8ELqUkj++AyAgJj6Bty8rSpcv5JEJgfOujXmtrIWKFcsptYOE14C+1Nq68+9sksnNZxNmI8p/
ovrtOCVL6wJrYCm3SiYvqnGx3Mkjhb/xvqj7XFjZxOJuS8EWBBr0bAkusSkQ4MXObik6vMzgPwbI
yNKn0Iavj9i8j/9pA+JiVE/rHjRlQwhswFGSDpazQuuDp7FsNTIap7FZMWfP/CrCON3RVfBFp3Fj
wmmHCPb/oOcy4LGhbskxCr+NBd7E9CFB4FNshQX1xhOyIB9aYfXgWDPTBvqpisWZkTqP5MTKFxPk
VSTtlJd9jn/5wsfL5ssVCMiOg1jSKvhYQY/YDzkBykWrOoBTygUZ8aaWGwIsc0RFWHA1FsBEvcqN
q8h39KPLOxppS6b3/uqdboCUZsW+UDyfqI8yk6LE1qYgpTTWRxCHxWpHRzp6kbZTp8jtIBmfHgMn
3e0ux06x+ByAzOBV2udBWi9QZJwkCIS4NqWbls2nhm4eE1wluGIP1ZAC5Mx68xLe3y7E27EY3RE9
KhpF9wfDR/UvC0ifL93O2w0iIMItlhfA0ZXZXYlXi/Qk4gcmCLAH1O63sDpbNs3qlvizCo71jO2A
jF5vJQdQLWo9C5xbdEiHo2tzzd0gX14Ov6Pr3l1r+z0zElOwuCFnQfuvHTR00cNpHBou/hMd2IA/
JbgJCENGddAphosgBMX8dwtFY+CKUcFm82X2YSgq656/zP9iMUswE0V0A7K/SSIVcWMh5CknIEdO
QnqTbhANjab/ZT8EwBADulaa149uwxWPVNivh6Yk2sQRD4QpK4PKiWQ74P6Szs3T3Nyo2qIOKWxX
lGOad4wmE6vPgY//Du3w80RxcdyVnn4sX7hNtN5g78r1C0w0y3Jo9yVjo6ctI96Hpr1klYB71h6A
nTPl7KCE8lwZFwGZERQY643Qas6Wlhb8C0tJiOKak5ueR7ug32AqJLW9Z+x3uBneuLbAqkNEnBiU
ubCvrJLh4Acv4LlpyJk74yTZKclKiFwJIzzjgFnLqbKnUnp/ijGIMJ+74MADR3oHCbEoXu44+N7A
0VVdTxjhMOKR9+xXx8JYnE9q4ZvS5a6c+A0Vnsalsnu6FCnAOGt/BWvJJ9Qv1cGxLZZLO2sh468t
0CLluloBfRJaX8UUblx4TKs9C8l1C2rLoXaXR8ZcoQ3Lhfj4MuRQJ4Bx1S60W+7uTSCJnTHRrO5J
CJuFxOm2kFqax64jkDN3n/6NmFzpGbQ9y4AClIXApMcS/L5EfP+UwLVl6lKwJrp2eo4J8gb2f0Xw
124wgZ2q6MeAcMM+dl2SN3JKSlO2lwpGpacS2IdRT6a488CfaHL/ChpB9+VU05EHdfrCGDDHB7YL
wMmb/S9x58mrctqIfvqECZDIEd7WFOZlNtQzzsRpAAp/ZhTkixQ4H1YnMhtJIEeDWVT6X3uHl01V
WmyWtjPpSfKRTovnDJ810l4uQkQqisf0FAj7Exz97+Ke6W/CksmvPFsIvvOwcutBgANIN2czrn/S
QrNkgbkfVi03/4ZU5tBVQVVPzub8iAee19BCAJmDiVlTMnVppEmjhSGChrml04sSZEuh+a9jxlWD
NwHkraVCLa9mJ4dEZKtEUn+0dPNAnbMA/q4IrYtMljOEajCafvR880uzAkmVtlBpZnRTSiYfUtGb
WXByIAh7PXkj9oD9q/Jss5kecPQYitBPZN+DGHs4EhWlBXepd36KBqneD1WK2b/b1IMdp8QvYyNl
0ziTDYwNY/bNAGHDoY3VCqehQ8LyOdDCBDK8prj42ZJRo3UMxKy+yk3D2PmrT6seRJMXdJjwILCF
i4j5h4xvPzQQ1zmMKPLQEB8nnM1LXH86QfIVY7ysGJUqb2KSfMRUtYvdrJF5GMjZacLjNOzNAHcw
H69Yo0Kg180gZY68VXClDPeKLeRUx8NJ1Auxk0jgRuEs7ejTsg9Y7O3AgUK5Gx826Q7j2oGA7/wh
kVyKGY47PlMJic/+aAGo0y81BaYPCEPkWDkwCkmLiaSxbxmuj35uL+A4/ujt1L9Idn0l5dXwZxtQ
UqzJ14N1ArBiaP1YEfSjyLYeVDNXEy+N2S4d/I7Lai7VLaiXrPRQlHT7iaucgUe99gbq+Kmz9MYL
p6P43hPVESzi+/CTOhtGSzzvtuzGzxAmztqG849aYnNYOegEnO2svGsI+wJaORET1cUtPLaYYW3M
5YL7rQ6rD6U/1oFGg99W2em4U7KYhcnNfxFKq62V05Cid7q0q9l2aqBQo8DGRa6KJmVhEiJxAtiz
jG70CNhPUjJ6ZZv2v6OBavH5RAmr2bMBh+b2BsVd4UujwuPbh0Px0dWpeo2SsUsDrLJbJ4vVIhtr
20cv7AE79zN9idVVQxQWHiWRHIjPFuSSW1O+JzzpBfrLxGBKoeoyCJvjN/D0plig3fD/WpN1Z4pQ
wljjgRITqjQWkJLR3u2qAA4qJqEmXPRCNMzE+OnQoVuDz2P0E/KOk5d9iaARgtHEtBBr+ejAorLJ
xRfWyneXw3LDhbW3+rF/ivzwg/qHIHMCcTycRBCt8YMwZPB97UrZFR9H5CudTtlpSwuGRWBITSus
RJ7O2nWmW62clkBPQqW08Uq4auAj3Dr9SKMmFX7DlyJv94Vko5Vd9HaQUUV6e542FuKk5XNGDvaJ
oeNjTt45ngT3VkIe7dXAUnkNJA/D6022Jfp8D/4xwoiFLUsM1yrN1q4sNPlBPu85qB2YQaz9oxQZ
rwX/bqlPLsd4WFHMiNw6yXLIjuw1QGgeiTVehIfubGQEIHNB2wmkv20vYdGYgi4U6pQWjW+7r+Vq
lzy7A6uvne3SiJ19h65KPC3WTxB6yKi86G6PA5+0BmuWZZZ1Cq4+VLAy/1a08kLgKCPMTYKXNMmr
ingze53/kYGlpKjexQ1IyM3EQVJZhYgNHL9vF8nfm3FsFaEG5m8tJslrPXEqUaEKliDq4nLVImCY
5LQkbYee3E+fOI0yIQzdVX8GKQ4jnaFM7FXDTGiBh4AkU/INN3gcSMBJXN83iAfEEseVSZxAnaWh
akYNklnTgjMljjQ6S4T/3UxVlR2xnmeYLJqDUb1l+qT1C9Zdm3QTIe4xC0HztYf+hd5x6pf7yP7f
CZQZkdkri4Y2++XkB5KTULc+xnPF4PGBKAyiXQd0srt8AAHJD29n4lTFoCAEq/URCDf+Pgbz5U6H
5vqruLd4D5lW5IKwlOVS0RsKDUIWBrnxY+YyU2zdDL26QGZ/6bjceKERezBSNqi9OlJQRysJp31U
I3bZAOoD2nlpSznR51YcKFd858p8bKv+2IYwA+81HatNZ0rvEQpjHlgLMfgTVsbTJ90EQvl557To
DjpMds3BrJBNy2+tDmSLxoZ9noQ11N2+DKv52rGMiLDvz5gxaidCMY9qj8dAgfs9nwvUHcv+deLn
M4HzAO6DV647hefjS1yV4hsQ7d4cKsNscc9+fmSdNVD9Ov2C62he4SSJrrXl7RzCjBJFD4mx3au5
AXD4KuXx0YzpPsP2qAo566I5NNmn5gRsZDuU9QhUHJkJkscJi2nn0EeFYIuJPAgdpK55aABDlCiO
xxwMJOxngOHd4iGtgTlVFEsVVDc38z0rMBZOtJfd4I2XfdtU8kI8ss0KFtyiKL3pRYXJmbAfbcnK
x4POtuPubFUDRPH5nfIq3NVlhZLnCj5MbTZ8u+mHGLo1/eLBkRDnDtBcKOkXo17Qg6LhP20NwH6j
HbAUf5+dtRJizB/fVVauprSXxNr5h4COEVZ9YPEyknPnDb1jciWBYAQxiibhJa0Ff5wzhGDNWJjs
rj+tOaAgUdrgDteN0PYtzKEMCRSJHN+1CVzctJDk6UrusZHLxebB8Ir+Aebvj2q4zlArXJ/aEURr
+ntasTGVS9Ky0SBQoUH7zWYT7qkJBB5uKtj6qaQfOnzOoyIxcqyumKPNCGorgy2zeg0kt5nRAgw6
bz2uD/yFT43syegAoxet6oioGA98G6AFoT0hO4hOFvxXNKKw6P2UGZJKxNHouHr2/lF0pcLDYsxR
gCT/+16MSUW4wx/fUfPhoP5U36wI6hdzm8JSCaN1H8Zo/nL0qfyfuVlz6LrmV2LMd8YIWYHFj4ch
DA96sl1rxdFKFK0geDUQziWS9LfkNWkTuyVZqaNJ2szocxOeIlaHZ9buAhLRCEvyhUUmf4aYcCt0
xGCwq0DDwhYLvHc3Zl0qd6H0SXex4t5gE5NCuUoeIFDKly/lk/rL7bZqMvVs/3x2qPfgj4vmDRAX
K+o1GwfNjNrXTyoGh1KK+tPnmO2QTM99dRDDkcDsOY91BfM5/iLDy12INPFjYy3F9mJYhcRMbc9Z
gzfoU5nh6P/0IpY4p2cDagyzWle/MsKr89sZETvmVVvJ5vHZ/kBlFA9ueiCqp4pnoIlM31naUixU
1tsIsZE0K0FfSi4Ia6nNHVOVxDziGiXMYxyc0wFnls0sJQg0Ce76WrEag3mAL3/8/iuumwRC04df
t4M1/domUytzk+v5t5KMeOM5JseGq5+LFjy9f0TGVoKnpjBhcB2LytfS0AYOJzmjjLRAzKm/4+OU
BsuOlTySfFS8pNYo8uKWkSoXAZoniSkJMEDmFDMebNYmtyb00QRKspvaW16Te422K6wbHi7W0UDd
kBkb9jv0ciSZtlHPl9PsFU8QOPRhOc7yLYHLwfHzGby/+pllvYDFUpfS1TNAD24BlQSqS7WMv+D0
9fQd58s0rmKG1ax4b2CkkgJPutAxJl5/mxvfIvNkCGXSUzFhMr51ECX6GcG9HmuvZ1LTcp5UXglp
zintFejs2EmI9DcaDA5+c5jJTvHgrYgO13b2aydzha1Ge7Gh4D/kx3nmvQO9Jnn4uVRcX5Icmjhv
0i0asCnv0Bnl8SDZfuWzedgHdmgz+ZnXwygRs0/WM938YNLmDGYuDgMod/cymMeEJwXvQqSWpAgi
naf2DWCfEWY9/rcUgycIf24xylGmhvTgvtpGnDZ6ayDpYWHgpTcY2LsfEHtdH1/jgI81F4F0kkFE
thdO5nly0RpWANw7a7qt3p2fHXfATgADn3xsUpdiG3GwT6YL5qkY0wIlCdfVcHJkhlePVO4cMBej
+5nFVghtpbVfP8ptRPzptGoccMf/cbA45H5lkZV//eED4tctLDTH1uPj5m7Oh7GE20KfL0FqcnI4
gSH8cOD32pyN81zFnrC+3MU8PInjrNcoyuR36xH+QdaHsrS0T49gv+F09lNAx+HGNOLjOMmoIdXR
V0HaoOlovx4IEYmUvY8f9icD3bz+uugH/NqqbpU+4yu05j7/WwruSC4v3+OW4kXWPpeokoS283Dz
npkPGPMBbDcsWQaT1IiQekQoLok4qEDvlDgIRVF0E3Fp0EAt9ryNuo54RExTWShXH59bmsjfuNoc
jNuK5R4TjW9v1gRJr9vqh1Kns6eLDSNMS+zPEIXNn5cl1hQYD8e+PSXU91SmIY/vN6Og9GE3szeF
/1BUi8iJh2NkflLTpZmVUgRvBfh9jmR8xED+iRoZOntZUuo4txanMcBQa07bDGHYsoD4W0n3JjZC
uIMsMUflQhenonmlTSLqX3NS0jOdH6I4HjNnSbiCpPCYJVctB647xb2ht/BF+XtjiK2foz7tEx60
AeCvCJAvJAc4JObvEHFy/0MXPMc6/nBvCs/w7MZlyS/Dq0Ps3rkz0G+P4fcIEBoCsXzoRRuKSBTb
GE7G8fEnTNKjSv70XkcmeGq16LgJmfYlk4n1anV0v1Jg+xO/22D7If4bhbYvaUTWmnX9QWNR+32g
JSPdlkDA09TyHDCMvqX1HK9aIyTl2hUBGnHoHng/MdTZof9OZShVrF9/DHrhSlPR2O/M0Q2ffIXD
kxpype4dA0k71+j6VmZyUJe+d1MvrNGSZVws3vWZIKzhZQJRGR0CXEDcd/OrmTXDHfIWBxvCiqBm
mptsyqvYZAnd8jhR4s1quqZByasVhfexegyMAN2a7mTAnfe1zW+Y/Tr/+IQVoKZTaU1Eq7s+GD8F
jVxhxe0RTEO9WG1zSVC0SkLUaUrOudv8b60bc26CEXxtuu/Ur3VEzp15OgrHDIpwTAssJguc021W
40tKcGpEyIGDnPGNSqU8aWp0sRtCVEMzL6f539HQ4j/GfxrrdSuQ4v9Vwy0YYcOdVRy6yK0b553T
6Nclk9BdlRzpUa8sZPbGK4RtpIMU2jmrwVgKgN6je00oCjZIPh46PpBjTOcqAzmxKyT3DC/TGNlJ
W5u9nRnHeBwLzgRBVb3Ut3wKvAebeLfnva/+NTbCxrdkg4IXlbWveELRSNz0CpJs7NKiC0ay5icO
frYKNdD+Zh1I74ZLMghuF637kQGn2tlumMis0UNf2xykw0bl4emr7k9SZ33N2/YcEY234otO6VGJ
/FKlbJkyMM652C/tGJ1drEjXZUHTLZRIvMwiCUep+5+knsHvOHnFma0dB8JvGZZ8hyfZgu++LO8v
3L014EjJFh8lyK5tiGAMPXgZpRRER5qRmE0GT1YCUStmi9aegO2k7BsKVMkJ83O++QYJsZwu4w3d
Za3Yc/Ij0QAPl3l+VtU2xvIj7NJujxGVEwneV8fgNnXZhrkD/xAdCFWObikXE/GsP2ixk27gVk2R
CEd5TxQlJpV96uHiizNjcR040jQtlQlQ19CWK8p+ZsiPYaqwMQ10OW8FQjveqDw7HmVEcZ+c125e
G4a9ghn/80pp/4xVcA+wF9OFYS/Wste3uS1z0lQgrN5ItXupBcXvwuWXa76m7yZ1eCfOPVfWlLU0
QY2Oi5h6Vk4ul7GNqHL5RhjcoTBKIpaAUofbIh01laK0fMpqAk8AIFdSGe59J6NJZhoW3crNr/H3
//zyNz/a/1JOlKADSBml2vDYZ0x53yItjNmLTU7tDVssgymaHwG6k97Ndi0Lsa0df8Uuo7BhDCnQ
c34yoBJB4qG+XEKELvcpnvUyPI4dhs1grOvb58rPGKOqLQMkPdTx1cTOzCq+3WDcPB2OJ+OltKy5
94qyJJbBgK1NwSVN6bxGpWZY3gi7qZGxIYOqQYPFlOmcapCDuLZyYbRyaWFoER24+YiVAwR21s46
FIkaeHy2+H1hgu+XqjcACG8M8VgPm5Vp5CSMahInA/YupYBkuJBjkOG/gMQhs1rbhBkWsNdKBjLa
Id5SeNW/E/SdTVRKHBGbbtDayD2ivV+0HVEhlPCPBEDeThwD52UW+4nRukMggK2ozrV9pHpjv2S4
ONm8OvQK8FqNMdlauxpiaMLNGwwOu3P5faOs202UazIwHXbkqKxVT4Z3MDVT5gUI1FQtSV36c7GH
0S1ySM0xVcKt1BGxbzf2LZZTTK/V3wjNUuw2nFUlfjI5Nngzo62cE3S8zN8dafCmFEJN6KrbScPc
Pp2efV3M645d41WJrFldZPW96cBFI9QCumkFfRdg11iapk/A3ZvMM0EjEUYBUCatfhKlK7DiTCaH
DhioJyYxONRczQSV3lhmXeUdy6jbzqQ8Biqz5tH6za64c8BdR7mfPa5xyPeJyd709+vppSWEK3tE
/UB96aHA+9jEcoFhfVuaLAV3+duPRRQHhZDBWDDGFlbSJX4vAeBC5tGbnnKKAFRQS6PdSO3kKLd1
QKICAVddIjajjRiWhYbRGS0kFXkEfvna+dF7l1FBDtcavQleAkBs7UcZcsI/vUSIl3/L49DY173x
6xgpQ9OmxbzcAtFnu6Lta8KWYguXeHmD9+HgsKeja1LhiZDSdWZS5Cl0lRG0WnVaJynqMjkgNa0v
tpZfPFb3MmrJXDJTp/3ZMK3l802OSDQySPmHERQCBue9l+niOTqpVoda7gYwlF6x4AofCYbid/EC
9AkOddC75FOt0md7Qy2JQc+kfBzeQoSooUJLc6RL8ElZjqxv+12Szxi0kgBb9C81JzxbDQg1bkWs
DWfBgVpc6BfVv96cI0xF+2RaYsOSMz2VPj5OAGpZSVfH1VtHXmE1Yz5dTxzz1VfqRJAP71mXiL+b
h3elfsLnDgYkEuNTV8LmpHrRcCt35gfwiUkrC8Sdpyt8mr4JTL+JIL7UGmBHZ7K/uNT9jHkHZJSB
Fls6l4VM4tA4L9s43hIfXfk1XdxJuldy1UqG+l8yqSWfZBApBorrJWVPGILt4truWuDvNZySLK/r
db9fcnLZ+DI6kKUtzRhVnLRceqt159aHlxxlM/zyyMklP6UQhGf5aMCNWBJv9F4phkMbCHzcpRGx
x+ccNH1snVU+z0uHJfTsLWOb0ObGsCWhu8607TTYuhhSs47/d/U3sL5ie4FepT0rZaNfVacJK00X
6mOHyoxSFKJ/oDkPQ8S1I5/WvYjDKux1eqO5WwEeMCnFKCdnTbbo1JGLAE5t/dtOQllomFLJU7Oh
wxsv0YEwgQUug+VGiLEPi/MQpE7rPlRVktZK72Hn4WRBHGqY5lc9RVKK8bxwK8EUQra+SsnO8iqJ
wn8Sg/ldmutvguZCSKuD1D/EhNZT8841g2M4gBXLu0Q5Qw13C1326DRoOv1087iD6ihYhwD/FTrh
uFJKfKWSFDhaCEBW2B7hKjjmLHEfmbDvB/JvO/FGB3KIpLx/R52tjTdVsZsUPmj98XQHeTLLFxgU
UQD5OPIwBo+G0hkAjltwTnlF1Swbd12ddfZOu8wpawWdwxo4jW/4sU+ZkaJNCLRUCZWIc/BGcxWO
Yk+FH05opbfeXfB+YrUCptqh8DTk0Yjt331ylvo8wZWP2sowB9tDSrOs9oZ3AJ2SHbG2qtzY15kh
sSjipcvau9xr8mftofhb6Ovjhqsan1IvHPiDAbWNKvd0GW8acbwHSYfiecYJKyS1/71f0qYujm54
gEeZ329Hllu+uQUd0sImrBBFKQlSxaAaeg/gJXKgxpCy74CtzHV8SA74nJKTxVv9c81W+SdjmsDQ
G1Je7bJdbOJ/Nme9r30SWHcJLZgXa782cIPgqGFCyIy3JwZgfk6XAesnvZGO9vptLvmym4gkxIn3
22V656fBFpgJeiW2SkYQkJiw9RUGqXDtHLTwPoNFa+JnYDe6/bGe3Ffvl+2gB2xpbLPuVIx8Dow9
+ZD4NZx2D0vEsAhqBRadyZHvpRZCyoBNN+RhAgL4JL2A+Zvedk3ySj66yk3I8iH6tboQWmMKYW29
5aJx2D7Gdbxvm+vGvHV2YQCokOlYGRbslo+ma2paetkUyjmBeRbaRIwOiM66miRbISQNneK9bBxk
fxz/V3tGNP32k+V44xjaFm6yK6lThqXfArqoS0vwEFMATyeRYcLIjo5VTBee+PbkwwNuQ+QTME3S
tv55v5zd1cnIih4trXv1tDa7NzEpDK5+pqJA5fOrHxuDxJQFf33IMUjXyXEZ++wu4NWRAOoO16bE
v73K1QzgzbDWwCmF9teI8RerOc1mIVGu+ASjVQFpvy7NmCLE9+/NCo53n34gzmhhUkDHIdjombHv
UhsUV0lcbWJh00uEJTbQHLtOiTcOCnwpwhIvGtHHBVPHf9/l8uL61TZJrw7tBFqQMDOi2hp/AjTj
ujnzWeJjfL68weu8jwdnf7+wjhrpPqrNIQ+BR/mQpRkXFo+Dh7uvQ4VPtkrU1fKFqBWzEPQTukfu
sJxjAVWlU8cT/GZOkS1FkFW8XfR9pOIiApLv8eo+tr1QKMbwEvH0gbvqc7McU0TvDyqRGbAH26Lr
tvfIWfGW7+cXVtUV83XkPBOHHTkAUZ44E2P13kD2JFuiIg+GBDn6baD1SXaSq2R4psTkIzklophm
AmqiFnNLp2PVnXFcTISCBlPUwpq5Zy9ci25fOD4Pjp1HxVMOHGd/iRExX84USUzaBohLWZeIIy3v
XouvyrkqAxJsjMapt0kyfgVyee9MV/TUQOmSRZtMWWCgRK1Gt1B0tzw17hVw5DfXqh9kRb8FrcbP
IImj/8dkk441hpQjh4juK0soFqrkfzYZ2rCSdV2zssGJMT8LAtWh27a+DcIhhiWT8Bq1oykEzqzM
Tld1mKLJybtM/iEEJb/Mh9jNjb68qKanUUAE0F1zFJmufV4zQCvSeRCd87mEtPJ969MEmsen5S5m
otOJZzEfmdaqM9+XQAdg6Bhu7aC2q+m3W8+gmYiqSDPasXB9QMgnQdhTfC2VkiOtNGRxHsxP2sn2
LeClkw5fYPBy8j649v9GLPSPez5tnl7UeZ5+/mpxsxyvrZmPMloXTWAFgVyZx9rEbi4AzUwXIt2v
AhhNZ+RLq1vtw9kudNIXHl9E3NFOgiunlTx8Lo+swq3yVxCrG7S9jCaxsRu1D+DbpfyvmDH3nMEJ
dMjf03/y3CXIrWZ/IqJAHi7GhV2QydXsVRuy7UxRrq26U2mTtACDcCiUNXYOTqcU+DeYzSySRfYI
8Pht9TmTWH4cLtd6d+lORQnypc9h7+XYUfdT9807O8oe6wNah1wwQxoQX3enpe6jQFdJy2bU5XQS
JiF2+eqz8idAbMvbJziZDYAPTIVTLxks1cGsbvtmsuyUvkiihj1Z54o8WsQRN2Qn96UEqUh4Lf/z
9TfNxJlDjDq1VqhlwE05GjlVzV2nT6uxPTpsMt9fyVAD2FzanrsP4SPZv62ATxP295/uHOK88WMP
QI8HUczlgjrt0IeBt1HwBgOGggwGzBgdrHuDhlG4JjavHu27TA33YivtCq+VUNwqtQXmat9tU4wW
spwYc8a3HP14JnAJcpxUUOrvUHHHqR3rjqtQqWbwtrnb7knuBfhcRpJ+sCuv21C1iNWXClKuRgxN
ar+qdtulYPU7NftmP7RlkZ0Gi37aWEd3UVLghprCFpcj3SWvAGjAHskQykf6gNF5WY5TAeL9O+EA
2Psilfd6wqvPYpsOC6FFaUeoRb5Z0P1EAvUbCBdu0IlcCNjd6m0uwLp7uc5hLwJLMJDhrMnwNplJ
sGtbUl+AtTV4PquaQQLTbtQS/t56SlJD+1zUH6R/rKnZG0uYXxSrPNW9Tam7xOsi5m6DgjAcj9dz
5I1iv8PRc+fnBJrHMhfJK44WfFgnc6aNmXg+KTU9HPuaSI4VN02ovxlYH8rMDc+765SosXdTSELv
b9zH8ddJzEKo9PEpvmCP5Qbw/VpM0sfGOj3n9foYiL78QEenxbOQt9Wc8zupv0byjxXf6Ld6ZeQT
LZ3Jcbji/RiLrYMU0gPnBUgbQXPS0uy3jcDNp0PBRqfaCQynwL+H1NRHaV2BDTgXwRz31dO2DtbJ
y1+9G/0obpVKvWw2oa7jCxDIPOaFIgPq2ulTpc4aOG8AGHR6WNWwgUH+Qgz/2EJT2klfoRZxEAwE
ypo9rWtjSNloPfx3ueQJHxCfQuyaPRmkrz/QO0Dld0beiR2e8+WkpxPMA9CryVVmaubRncMHDN9c
2cOEyNVTLcM0Bfg3NBPmUphM9R9h9GHElzhWjW0SZxAaLoGyMM69a4V1TqEnpX5ktcW/pWtguVJx
oHf7TBeTPmXOEFDag3hOsZyTJcjvXIhmSFHUtPntF+k+Nr84pn9w2VoFiNGbWSelTip38EfGaxWO
mNasyV5sTpecvVDTz6xO7/uhLvLaM0ApBsdcNdhuJLpMex1ONZEB4Qn3EITpMir7c+EuZDAJG2gn
6q2b5xZsOlwZw0McOkj4sAVVnYR41d8syJe03RaDGbPciWevXZTO2knE0cu3KLaGb5eJYsrS+XWH
V85as+bhvRZoo0whoO8WPC0XrwFqT2s5/TY324CjsPQUYmRW6pOx3C8cfJvJ602SjmUiLMoN8Ab2
xQcwDEo8AG71zFb7Y9EYz/kKOPs4VH4Uun6S0QzBDcCcMrrhtjQySGteI1pV2R6JOzTnvNoP9sHe
CoutFdv2U9TLhw6ef08wJ3pQh4986SjUvSPP3dS90DZS6pQCblz8kjIQIgFIc2tloA0jvmdF3mOl
A5g6uoH6E8IchISN7w/Rar+WUtpBbg5f+hugmbe014SaA/Hxp2Q4OQdB1+8Mv+cAQj6WzMv/e0mf
QtFNp9tgCWC2UjjNBCJDR2bMRysu2JVeSPra/5vCudzAnbv4tMwN9YQjWbneE55xpoU0LaAV+lry
03MH3CvD586y0zPZJVZfEhc/jxpcXq8lSZBbUnwb4jWMcJB1a5aLp2YICX53Yxa/5vF1uC59/M0Q
QIGWCuAGoYf81e+Ycddc4uEo74+tQX51KkJzxJosVYjptWyuR2Gpb9IZRjd1H4TV5t0UZ61D8p0W
ZewknhhU0YcAvYTyCifRlhjcRYPZI/tV+4vNAcoLr3erBIbWPWf1iP81isLx/2hUULfR7yX2iy8k
s+5FDQGNx+8E74FjE0WOFytY8oFy8S3Vc87eEOv7UtO5ymAMJPswP4kNKSahaZ/6ntb11LIgmDoU
Mm4cV/b/JvJTaHLOPMYYROLOqlzMcL87Uvm8ArjuAHNbvKfIb+pwlpXuyAunpiyFQjDlVPv83HGm
goqQzIcoMspm09U9rrNm/eDcxRU7TfDmdDVGPgb1a0kDjPn5mipdSnNBHEFRa98AhQ6LYJ/M+oAx
jsoZWtZab5uaKPwTLMElQ/j+t8zcODXHg8nE4g1Q+T7Atg2Dnc4/5rEm+euMPhXZ7oWknSvI+gwU
IxzKs4tpEIEN0CpX5Oi2HJ5HJ36MdORZdfqjxjFWeQJH6K+tTOH00FrDKnGKY9z3Y5aXOHGLmTOm
ec5OZfDRDBnWJ8e9JqM0dAMLdx1m4IUOiI49evKxsGNwIwUSmfXtqIkI2klrDFX3Z/rs5ohgswhs
fnPELOcfSx5b/bUlWbIHwrSMM8yQMFi1iqmR0WBdXSZW/BWv486bBLq2U7Ce7raUuc+pmkzbi1xE
0JZ+eaZ5F7/KOZXsPjdouURG0+Ueq41QPHOGlUpKGPXZAyXoic6qwp8rKJkoa99s0UmrvIgdGMOR
HTy3GQcwkiuNPNKSPb/rbRmLciHsVRhhKB9nqlfh4CEE1WmTEHr0N6tqQ1s/74CTWWUrOLndkf7Q
1cQG7+vYEPK7Uuwykw5hLkKNfVK9fjGn/uVGBXKdOjRKYVJlgabK8/taNyX57KAtsmq0Q8JcSmc2
m0Y3ipn5zOCxiHfj+tTvSKzLD1eNMBN90eahexxWaJRK/vXrmuYmUF+5LagpnpqVCle/3TNQgFjU
phnRr1NUW2s1cq7Z6Pcmilhltf1BJYpUwjLZCek0byUFrOWPc4NHwyLzLi2eOEaA2NU1oQC9Ot2t
kwBSKW5HJ8/j7ONKW6acCev1UiiBHQsssGnXwvG4M9/FaO5jutJwrf10aStRrWls6XlkBjsOsnnN
EJYK1ZMpcPvseO+bj2DqU8Johp9woX43mRzRmwyw6m4RtYAzyAjdJWJ9iv7eeYXmTaU2KN6A3Euo
eXR1b8pr1HO1a1f7O8XezSYeFbMBFw0F0cwORlX8etvHzSPcKCbqT8lFIH5opCbOH62vbTUuQbVU
xSMoxMwwYK2HPTXo0ZeBv1Izuf9PbCLAokYqa47Oy7O5E3N/zgAKr52DFamqEGjAaYyBrcwvWPDw
p7uARi6rsBTyovz9ZkP6sYG3PGJAWzm8XtHZoU73ZN/LVLtgFWAZWiN9BPWaipY5kOoRnvlYsvtY
IVRsdKy1JF0SnOckMV/e0S5wLCuMoSRHDqaxJg3Vd2WhtmyUrFWhITAeE71DINoy3vBolOikjCve
azDLviBwlWsVBDef6eM1+7SJqGpFmWPWPObt0WVPr6QahTBpdF0B2uNziq8hE/m0beuyGxwApNnq
2Qu7NkpzKpGOasIpKY/L8PC5yvWUBGzYfccyQASlSeju7OX4OxDB0e6iBW39MQKuqpwg4l+WXGcE
91XsJd/VZwzrplQOVEXG3eXMgeCSdXJ3sS5ghlfKx0nQjuqLswf+M4qhkZA/G50sNInbzfbedmd0
i396b2HzPMiMgFA4XsuGjJwYuN5hqBN82MLpiLrGDkqql7xwjsop0eTtZfToGqTBeL8SLPRsDRtz
JUGAPElwS1OyFaMBVvewF4SMbpt35OjSMT4o2a/Yu/8FDMhQu37dzbCEkbzz4uKheOquFVTFqHST
p8PWUr/BrXMagiG50iTtbas+jEXVnOhhxBq35ZKZulAmIR5/HCraK72luePmRIjHTJ8SzqGm+hs4
4WXKIGUaHTNdj6t7uT5DiCzf9PGQszbVd8t72spnNuV5u3LR6baRFLW20hdUrHrXnkdLFgtdjUxt
NsC6K53DLvqKOBtsj4oV+HSVBiQZwdmGZB3hOPL3ML3ltR31xT27s29e73UDu0h9koMlm1/OEgPw
WddueI8AP0BfdmFeXDv/Get4jnQ+esTQgOeKTgNtNjtaHrW3jZ4bFYm+vjS8Z8k/gin/Kl+CBzBc
SfLUlvOreu10g4nrH7O4IzqDwwJ1YtrDpSKBUbPb7RMyufo+nAvzfQMZRy9m8WzNZkoRdInJi0hT
HkNKWVYvC6UuWi8TPjo50r+1i28/f+vgC4K+1pEgammwogCQkEEch6el7RruQbLBJPa+yvx2pkum
mJRjn4tJSvkDjc1IBBZPADN0g+1+2r4VWXf3DJ0w2P5NFvMHQXYGULg2xT0KmEumoNojONMcSmzJ
QHYgwj9tDt3qI5gCt6zz+mPo0qPyUEfszd722rSKfNZaKq/YDvQKanxgOF2RFo4//+7OUZImUO+y
vjOpWv+lW+SbCLYHieGsUhZYodCrQMA/PveFEr0stPh5y63klOnib3YhlmuemOy3FqmBOLv4/fGa
YTPYrgyVkDq4NtXrGx02auIgj/ol+ibffBxz6l8ccAiWvUUNRyn4wMBWrCJM+pmjZHlgf3u7OUse
Kk3+/TzJHeNGy8mAagYSGQfFAX/sKKXU+XDsqZzK0orarF4UFeNDaO+81diYU18cDlZ0SPUfe+7g
jSaJYfDAjqWzZPzlrb8LzTuCeQqF3nb+8sJbT1oEJ1mvV2CLjeIJ7H5/4D7aiLczly4s2qoc0mZR
chjJih9k55qOK3Yp4GpcAGXLGQeYsi9PvzjspAKQuQi/iL6R1c8DNSefjTWZE+xoxq2KyizBHuMp
Tebv+fO/KI+K04YMh7mwpMUO54F6LPOAv4lVeP/+BN9zyt/oyVgVU6a135aAPctvPj63ar+sgwqc
TGaZQu+rVA81r/YTl3icKshmvI4jM9KMSgpUDkAH2qqSWDkJuwkthiOC3uW0kBQi3N/VP7fEslKd
0V5Ar41rXVZl/IS71Mm1ZDynge+xEFrc26ptif6RxLRmmgY94Ss8T5Y485CSSCll3wXKqmzm6cRV
ykMc6AKEl4c6C9j9IoAuu8sQQPV1/1bgxoe34ehC7nyUUB0jcI2Fg+U29PkbQz3CRLNvDKWsOVE8
Bd8B1z7keG+GrvGwipP3ZbNEO67aiSXJRSW+//QuQHkgSFqeu1JDgjdQdYM3XyekkmjAr74UlFc+
s4Kgg/aWWjJ/Hx2MYaAzn5xkvtqopsBE/8e87bEr5zUofizUdrrDX4HiTZGxxpiNrDBneLLd/YlB
gyRNLjyrrZeGJO+EIZkNBDNR7WnBOse8Qg3jpQQTmzljbXucAFixb8DqqFtaO1n/AECmmzakDYgk
RbExejehidHUnlVhSrxZy1goXkOXqfm+mLvsAvvFkyETqUtx+d4uoKpaYhoTO+/9z8htZc4Jmgj4
fZFGTP+va1VSGjrcYue2AVenYfGkVxQuzbSpYifBgb87SEi/WrKv8Hg+0Ds+W8xyrD+Xt5F6miJW
2OSdQbEF090EDtdYDnYFZdNVIgAQu6wdWN4+FS/bWU74CEmluwsntbDAxxONqdZjNJGnjHB1IgvR
jXJvZvvef/JcJTby6Z7hLN1+cl3ReViKAH2clX2VWJx8Cn5dcJ19mtcgIA3RH1QuSq2+SAN6/qdn
unf1l53IKxp9Z2mbEw5kn+PVyiJo1vcknn5R8RMBj+Uw+yb7LJzRIpEZTr/3P6xc5OFP03YcF+dv
3awZovqULAp73qZzgb+9w36IDzT3Ng6437vu5m2ggQfzw5C0bOQYebIqY9htu0zGVlY0+LXpx/iV
CDj2cWUwuOAsPrT6Ah003a9lOHSSGeq4uUt8bgDOga2iNBCLYCImtyCcVwM7XwfOtOetrnu8Gxas
+6yqlf2D6kddswCCUcOxhYYHAp+NXg9F4M4gSNV7xdGaOEMp/2JVINHN12gye3J3X4+Vh+6eqSaT
H5H+3r+ZVqt8lxBU9eG50LcER4Wl7I+lqIyALkGhRj3Tq1513O4PPKTIh8kOuHxziqQkT5UMok4N
QLQByfdoJLqzeI/gDWmOKBaHi2FohKaORpD9njJBbFlbV65c7YzUyVkJpAxbCf6tV7DAQVW5EB3Y
PXjkHSpo0MUormte676iI+bRpBoGtoflbu4rkKlJTNo2EsrkbcOxUxXFWcsSD8Gn3e0pmjNS1PyD
KXOuxmzII2Qmk+v+cOz0DOvs7gEGEzcHoz3DqrL/ibf0yk3NwAeBm8VAbNEZ4WaTja41hxE0fAFr
ugTh3MjtJIQ7OopTifa2yqOyFrE1KRYzzh8n00AzSD3OMWoo14FCOKGsJMBO8iDSr5FevNQDr1is
GvP5FLNBM+Rzr7+qMSIbWPxZ7skuplnc+cDidsjKbkubeHZQJm9tQFhTm4xXwZeCtn+7egFp4fKb
LYnDYS7eC9E8oKAAydy/cePvjsN10V0nbopen0h7XQCgpxyj2O5uNSlLTw1HwPlmR0tLiuxTwrVK
3FupEit2InAVbRFapPgGbBlaPwHtOV/5uYuJ1uUgCgczRFsKdhKxIwsBDqfnPzw9L4qAvVcQLv/u
YmnwlIEg2vL11BHluiIdSNUW5wZiC9CAnSl9JiesoAOtr/gA2LcwaKklEXyzRfK4waj3jTxiqNQq
sK6jwnaja4LaHxPwrh+KDTr9sG8RDtjtchWDxw/ZGfBC+zpigNOCILqSJmsaINWJyZdN34aAsEEu
yVd03RV2wd1kbZtRkvRXXdKpafItiSFmsq77qC+TRj7k3EEotdM5WYYkpC22vYH3kcgkwZqMG+5y
21mpJK1ezzBC+MqJOxJ7yF8rIPkjXM5dm4GF7dGvrqlg7TP3DzQfLbuH6p/HZRY6eWC+JItrgWRe
mDbOXlgRAmLiEUmmYf36m2wyGrn6azIzc3OiDwLfGqEi0A/zLbHRu9tDQGdlMUSofefbSnSaKpvA
BsSTPsN0PkI74OS8ZQSv6baSY+ex/B/ptGy9CnXmxD/3dihzEgA7rIRW4x264xb6/Csjuv+Rfndn
yzPmgMLKDna9/jGGyTpTRWPqaY/hvLFT3cD8cM3Xj2SYOUtgpZx8D3y6/GHhfeCFcvNoU1Jw+UCT
/duEJLoa2Iajhaim+XVshdnTwmm1C1EoboUsod2LgejyYBe8qx06l2veZV+KeF3sGU5JGXCoP2wG
UJg3UahMnoyFp0wxkexQmxWoAlg71/Dzh8U691yPf39hSRCONRyaIBoIHIqnSr6/P7V1cSqywbne
H4/JnerByxYQzp8qZJRJqimhNTB48bFdxcPorYdVbGEksDaTDHhR7tCyovb1S7G7LtFCvlg5ciRN
b55FWU9ACkb7mq0TwwWonbUg7r8QqY2Kd8Y4YM1Hma67Q8sYQ9jp5MZcakkRk29OWuoCoSuMJ4cM
49RgeFc+IfCndQr70nqJ3onTkJG6/54/oigo9bhUnJgb9bmEbi+sYXIHsi4NBe8yrvMtAvUajUa6
KSEoeWcs5NPmhn2g7gBWQO7P/q9G04puScIJKZiJ4tq41wQyUVH60mjAJNa3uvHD/BkcnvQ2S8HQ
DMpy2NQBob2MuxoNlw3YlAD5ZaP9ShFh4ZhaiupzPr7/HIkrciI26MxcssdNF7DkbWxAAaIJENsw
92mbJr5TgEwUWf0icq7nWatL40D1s6+rRXnzq6zunXqtOmf6Q+bihFNrDVAs2uxci32yRhzPrr0q
5Abg/Cjg3XS8OV5VMdWxLGvUAzVmzWEm1UckjDKwAgvHFtKGg3/f1kYKHzgDA3uXSMnImNo9HPIt
VCHOALIJZWiMG76bZI0esTxaiehSOzqwFBNCvsdMpCSfwC5NSUH0Up76RnjyG9o5Nz+BuWKKsbEz
9GULlIT8A9KtvFw/VqrpY3dZZyaJdj2B/26qEoI7SQ6uTwZatKQ8CBFzytWWP1WisBp7FQf0wsqx
FCXF1T7jMsgkYbpd6RDjVq2FS6hZIVitgA9pz/OjIf7HYpHlPbKqGC7b5ByPOL7uEu6TOqHvoOg7
JYJNG5/JfDJ/Hc8ZLSnhBNsW5fUvdqwcpOkh78FtI70NTozEkLFrEG8d8wEr4qcIYPccc4skd7pQ
LjHo3ihzV89c9vti757cdohPJRmvMih2juKr41C6mZ9XV243L8HTAc1jmVPa/uzOrJxN0R/APDA7
k6EHFnuNG1JufeApaAua8G05SCpbKyYt1IOUGiLVukawLlLBjG/+qSXj5QbdLAiOnt5W4zbETYVE
ue/NfEmrYMqj8Gy890Ke/NY0jU+Lai8g5up7/38W75SfBWTQ+YW1GSVQjOb9W+0DAu3/F1urBb2D
7CohRwTvHNIJrP8x2QFCSVLmLWzEXF16wzcU7hT7lAqmbxGVLrzjcv2JbeBPZKqtIBYsUD42kr0c
7eQyHGxaVFXB36hs8KNjVix3irGldzCgkI2s3yNBYgE1ZpEVfnrcpytzqezMK/ZC0mGOesS3/OIf
Tcv4E03zDlelprZR0QpcpPfG2TKDVlfc/JzFSP3+bAMSXBcnRu3S5rLTQt6PJhHbsdXRQw/vuO6K
Ns9yOS1lCcbLLPrL1nskIePpvYfaOjub47a8zvtJ6d5E1QphUcpe4HHw8Aj1jy4N6mB3SI+LUCWJ
HxVbNv2VPdWW7aOFeEhpdYc+Hq5exB4ddA3ks5cW/N3Gi/B1P4GHedSL3ILZRQ2Utl5PcZD/mdvB
MtR/dNvIGVmtI50YC3MZFksppD5EtmYcY95yCljecYhh9phamUCVL2M893Yfqs0etGggieDJoZGL
hrEx0oYYQX/UmjVtjTk/oFtOLvl9TYX2yy6gfMww2KBc2Mthe8odkDQj54sUNR6r4lAoeORIyI1J
G6Yq1lGEaFXCDgPys6Fy/uDmqDOjaiGn5UDKvbwX7IV27fd8nurEFeDn8LB+rP2bYFTLcxofGSL0
Fv1M4tFTQGMqI13YOVFLpFs/WFCcl7tDDSaEtpURASfjM3fJNVhaUdXLC55DQ3SrwWmlM8X+iBXv
bcs382CDBlepGO87kKqF31pFBSt9gGcTpdajqO0SPN9baI6I2p/0TXC+M9tNQSr/Cf3ylvcI2kfO
dSSIfn8+YFM0URRbEN7pQApPLBDPOJx24mvOBkFhq3B6dRigiYOVOiLLtog3wMkGEr0ZJOHjHez8
XWaDrbqwW632CnC5p5O+ZjpYxm7oUzPck/hs6K+o1dBnZw/AP1pehfwQ5AWkvSwcXvPsWOgBdjdE
sp2TUri0FeM1Xlj8B3ka7whasuZ9lEE98pY0Q6l2tVH5udVGPyY3MqcEUv5zQXxrYYx3xAz557Xd
/3GyZila98jiISncTSm3RbmtMei6j/WD+WlhJU7ON60/PBsCfVfvi/hCa0avhXiO/nJcYtFLbklY
Xt5HIw1Jt0NOKv8YjCp/Ed5ewIQdgcLtYrn4vyh1L5H50F9qQTppoDH1zlcoSj2qVSmcLufJRXiz
PQy6TgLic4Iejs/PfbnxQnDePmWGDakVsbAd9vGODr/csRlZKFo+MPYHjjqE1yr/fUq1IFc9MlSf
KuCy3J+cxmW68y2AzL/Mqn+vN+TxMiU++mcbwpsAcqq+MC+/G+7NB3Xj++Qq/6p5K1lu3Atk8NYJ
kfwJXQZ+R4YKLc6qthvWL6uZVQJfHhWcpbZb5E5dtJLYdA1EzjplfZ8mBooy0uoLTBefKMXMOYxS
0zUNLAl74dhPBHesyXjJNjsf1YMqtEemREY5k8mJ3fdoZDmFgssj+WtoNsJfG9R+TFt2gHhtHXi2
DphbqjX1Gd//KJNYUjZOIg8iVw1c1XQJxvLNawVmGg9JYnCzdHQ4rNUNvtcseMdIFJivHNtGH8Lg
E3f608M+nKBhMS3S3roqGRfrxcT/7QUzBcpjuJ218MKLnIeMT8H8awFmzV7DBgbWw39VA7Ynk8/f
H0Qo7K4iUqffLHxDtL7OoQMDghGGXyy58SBZ9Gy0CKBhXNisfxH5zdIsUCxfAQD14CdD0A/A32dD
3f1LwgPYGo6owIU8zZsrn+HyaRPtv+vbceTutddvzWjrhpfbqN+5oVmXEQX2h/xh2Xt5zAl1R7MH
NWs5r6XikX+TuCd12yFCGyUS5BCHKDJK0hIWXVnVp4J2oeQBpujsahnha2HQ7Zp2BN8cxJf7DCeg
5m0nu5cFbHmfjbywekHHCGbOT8uBefm23KpKxOezcIdg92kqLaWtgqIBYg1Xf1MMQu6hTUeoM6OM
CEjMg1hErxS8G9xuAL7hDo0rAHuY9CezSgpudrlc5zp31F1WA+qrkZutQSZavmHYn8VgbY6eq0Xx
mZq5u0Jq45GgkEPtKx1fKsALWS5D60pvZhaLk0L2gmqFAUzagBMnQDVfuq5/Jn28eJwjMnPNovOc
7tGJW/u5PxzshNjnDLKe4XgOYbzjz9w/aDpG21AizoDixmsGXfY+FgCCpB2wVZGBBZDtg3CXVKzT
zMjs71JqGNLMOrKjGP+GkX7f1vwRYzofLQdNNyK8yM12BeveOVrCelTBhjfUiKmXKTWIm5CB+HMK
XsYxKVVy4Bhy3+HHoj1vYgaJF/VI8BcAiIXnp4Tnln+ltJYyulCRWoVQNft8wkJjlVovdL4x8C8U
74bA2w7Aq2/+Mguo8z1itCWlnJadjcMdYRvW8D8LojcoHJSoBFaqACEwX4fYTrivKmCuz/79PmqL
Vh8IqqW/vl/FF8tIlmV5QnlSKH4Trv/hqU9hYQo7qQ8X7J8vwmnh7dENusCKSFBhfEVyA6oBENPU
3HdEJ4S31+U8lKUZo71g+QW/ip5K/YU8TYn+LPtbzrJy4ak5BYXVY+MYRK7ndVlwciBGaMF3EoNH
6c1AHR5l1iztnIc84qY54JjyZE/LPPebx/rSWgC2GL8r+tgFspOVUs74Y6dwdpu3BPw4xlYIsGqb
anoAIWgbcB9o6dzBr0Oxl0R/aWuI/Ey7CdTTVITTDR12ilM9S+em+f+SLtUZ1aLyGrbiwA6QSHH4
VEl8eYazLG3lfRx4MwbwPm1I4zQnyEG1M7VwvNCdUKVux4+0KLreJPUxq3g+r2na79X3dwK62qfw
X2uQG/Wva5j9/JWv7NbIlmzxEw1qGMTBJCuhsb8EIpu3p2/gP/8kMOx8G3xtbiwQk4GHFSo9I3lB
YaHVurxTwPhmpvPIHJ5aRQ8SItacumFhDC1zG6ojY6T+34klicxGmVl04GY5rICTN/s9JY3tQCL1
dlcCru9fh2yR6TWMhYCDBZXoFG4t2DD2sibcZIOSGH/Gb/l5ItWYBB0SEO1e3ZSZ2ia8qf9a9LFQ
GM4rtW2HkwdNOpW38TBCL8rjP1WnjfT87UdVU4vuSH+kUc/aB2Ve/xA3e6ZYvTtteplz+ZVQs1SK
m5s0vmLwa9Ep5asEgxh3pO2LnS1b5N6G7knPb3V1HSfPe2/a2un4u+iJtvN6I3O55AV+jEUSttGs
SjqBxYuIobcGwOso2VZ4d8/TQpw2iO+Na98rUB1Q4dQLrNkNA8DfiI3sl/zHz50uPKvRH+IFV0wa
1cEAXxdyXr85fPLP31MxGyd3kfxiNGlZCCZyrmsdPibWYNzaihOvCKIDbsCAa3x0uCspsvCiOQg0
tA2WUD9fa+xSoXLUatk3x+BuevcKwoHMzoo03LbQlvamF0HIEsqeKRN8fml54vXUdccG2tyjuBYf
IW4Nfxa6DzfZmDK14RBJb1rQA1LdSRGbHnN+/k1qx1HY3fRv41O3TWxy5p0UyYdkseqCWNRtfbqX
+7RnuLrQBLP9WzTemwDod3cbzXgb6HuEd526g0/LB9T5xOOK7TzZCdPqoxQpvlgxZosls09hyXAM
tVM0G8w9tb05DHt1mPUkt2y3M/DC2XLDnQufkKjBpdlG+O+GuwLYuL98umJ9/RA4HQsMaH+p9lKO
IoW+aOgfWrssewhyxm6ww3n8U9fBJgaVHl9BaFUU/C9UxFUltMVSMfwDnyva6N68SoQeao8eYW3v
Oms36En262JOnXTJIn9JYvvBD3y1hBHyiRu3IlTdFcB0UdaFgWYIufs4lErNx3XB79wvow7a9fwb
Fy48FZhAnNvdjw9Wz2g1EeF2L9G00oQFnu4WvtZ6OCbsw7aBJFECH6I6vm1oOyRT3cKUeNTBm34K
HJQBZpUTMVdhx3j1ws8ATvLYrNWjnNtKSCQ6nT9uCX4a3mj3AGF1CumNqrwD5lNb9MyVdCEXKhmc
2olew4r3JUBjg7dFgrxXENzsQFo1s5e5zM5+hq1Ax6Yz49JjGUoHeKHDZsJ69FUk3DxQOivCTbEL
d4Gf3fdFRAX7TZvOTK0q5NjgIQ5YcfZ+nzI5pti7Ke5hxvpdwXaA+gqciIV7pI/UPc1bKiQkV3Ne
CAVXNzcZD4Gh8ZCOm+b9eLmuBdPF5gpuYH9rirYrRmk/EmGAP1pP+LtIgtBw1jNrV9oPVe/FNlkJ
+b5wDvY/HbPHldJ9MjdEcycr5fm35cf+q+yPgRzMka+kUURocwUp4GgTDfxxl1GmaxINXJL5SLRP
cYjcw+y2A/c8mWQpxmWYJoe6ajV/xx8BWfQldD961Yoy/k+r71ytmeJhZOJkVXQU8D32M+8Wjucg
ZIx2qIoMElGIjqTMKQtMhOGHsf9WoVm7CBUiCIfxDyEOgW+qNL/mDirW+tcuWhk7ErJ17QCSb60k
cUj/BdfqpuvDOY3x6LDL7vNheaySyzm/LmAl5ZIKz8R4wZlaESO6+CjBR/f6IAo8eQawwZVawMBK
rDkgH13xWJHlXQeBf14/U7j0JyTmw5cpfAs4zDwHir7xH5RNWzRgmYv7KDH+wefcXA/UibqDBnsp
CrwjYMtxr27kOe/e7ulz8TbcrX1n5aWs4tcnEq08JV1rqV1fO6ajUTE3s3ttHQzGinJNbOG20/W1
7Qr1OVIboBadXIMdwCCAWLZoRk9FB/l+YfIGIznzNwrzalWoF1snQ507mQ60HW+KDtRCUQUt9kMi
dxAT2px01JhrgOdNGwxsH+MweihSE1i6AbDIqU5Cc/KtO/ErXRsf8vT5WD+Ig9B/LJiL6KOjSaTo
S6eDP8ed35Y/HNYhTAwA7QcuE76pyiWUO04fNKW7qm9rwpzNrlCmyLOmQNx0bLyxmA08HvOaMID+
Ms5HwBYDO2d8b2zFJKE7J/+NClxeakE0lAKCUPmV9dqrs9SGBgI+v2FwLjPvQ6K12ArVN2hrutNq
hxxQ5d9IKRXz9dCUK1f6NSpR/iyXQnQipTLj+utS5fnMV2UKOOjz+81i+kAS4bqOZh9+dlts4A/y
/BNEL50zZxsZ27FSSdvlYN99AhFg5zSyzN5J4g/QDuk/ulZ9hQ0rllZMiRL1e5C9c37xXqkCPRYM
CHBTo9V5DL2fcUfv4aHZCOCwMd+RygrJkAyxgkb71un0jYMXKjrVdn7h9RKTW1+S6/Y4LiVxJkJI
kxfp4iEYWd7Y4CRjqHPn54u0C9mQbbdMWwQjr5W2fDIgkKYg29BbQB4LBa/v9LpkxBmur/xv7c5k
yvzGNREX/gOkn8P5mt4uEB41pf9QyJ3/NhnSKxkTAg2Ht+h9hJtvkpY9jhUN0/MNjYPppn/17DGG
hHtJ/0aZL9CYMUe8IbWPo3bh9PjeYd5qrtHhUyrCiRhvIf4CVEnrQxyBtmj4moK142jZMG0yL2Iu
z9ftPuskl24evp2k8x02bYAozYeCgJ9iAfXflQlWLvL5JoU7w4FcuY/pr2QWyHl4LcSWziC7rjQH
0tiPzJEdqT+TuT17wNyemel0APOgvicfJC51hkSj/dtaN2KRc4FQuqNlfaA0HTABxOGa7GYzXKbq
MEB16NUD5v6Sr+/5elqgBAJtPGnRVKsZQztsX9HM+S69XoP09K9l6ViBLeYk8DJMDEdA/2bk9bBW
xPkrzaYkZUPJac594cU6ph7cCpB6RTC7P3LZ/E7E9wJf5qnBIMoGP6DX1ygv2Q2Q9vkRK3YiAzxe
hVgSyypGQeMNNlA1XyGRW+zf4PrPPgQgwbVI4BzRP4volyhyXe/eAWUy/BHlvmFXF8+vMuiwhYEG
7q/nRR9MxpjcAYTPEMPi5FbA2Klw4lVNElw/fI1wTrV9v9KcY3tBXxgVJJXDzXeU6feAUjh5IbYk
ylt7BYO1lpOGHK9y/fd1uWjlIqQsHPfjtry6xyPeZs3MIVb348+HVc6aTRUS8Q1fRtkmW7hVn/mf
5fgWI6KtafAOPQZ5M+Nnp2rPgBTkbgYd/HJ9ZpxSvcPVa/Kexlr+kTzd5PhE98rrTDcwWRKn//2Q
lSPBtj616pw/gg8xYmPNwBSoz7lDUSjCuqlXKUE/5zIc9fhA2wykrcgjdKUT/4TsZidn68FfSjy5
wsbwn00WmBEn+oc7cADF0UNuHqtm/Sg3oIi8/29v6HoSgbAYnqGoGuzq5u2BlKissI0nmAIBZsY2
yfdFEFNVf5j1oSpHEQ3/djCRfD6A7Umk4gd0psT0BqRk+BiRduyhNu2jozmBEngPPA4WhzvRB+m5
BNFUhun5AID+Wmbm4/M+6JxQInZjwa4CwdzW+9Wu64oDvJHvW+MkmJbBezrlZf2Xt9WkERIBcYNr
jP+wR2sH2EpYLZiEdZLmb9/nGX7NwLe/UdWrjKmvmrVMErDVjdoP+E2WPasVgtOGr8XzS9esIsKK
xqjmqp9Lhb/rrJaHFUrN8fgQ6j1dFsTsH4P0KrjjMqmqx+Nqstxpod+VikIvcexmjXjIQYPVXPp8
RRrKwEGtM3fEPtC90Y5XBF6Ufpk2ULweEaW93qVFQG7YW2184l2rjhL5PfYRfRqfcg+ZeymuEPMz
pKFkQyRldkk1iOJfMHKCkWABCuhG0JIjEQjYp1O3adax0I/g/3YGpXvShEUEPqZ5iqgLOkRZ4kVl
r/PsxsttAdEVoe6xIYBefHBqAjMkW8ZrnuWv0zf8Hz3FEVhYxpaS4kOJbGzICtaWvKzRh6zbKv1z
mE5h6bAPyUzhoCFSFNmxYs0aTVVaHqur39sy+L54CNj2oCW2tff94RZXhlzfuAehm/xRjgJfKvk2
B6pX7EFQqO9K4dOPhajo7gwbXDmVMM+Tcm91pS849DqHljc826bbnDinKIi3boKFEeb0AryMlPEZ
/SQak8gjG73EhgZ0Ay4CAPGrAQznP6/Dt4ez/YYFRFtx2po2ITvwVxMsscy6iwslE0flZNbsiW6G
UiV5wefLjj2dfSwUXx5CcavK+dAGAWP8bnwB3aZuDKAL+gEj6StMy/qbpE9PgzngfGYBgGV19H9A
c0NpxrYRd2P0CJLW6prY/oiHCLKLYb3+fT7qpxofWMZa64xd5htZOU8LPzhdOoBKVnpurA+5Fwo8
MNSzF1/G9yJz4Wleue2TxBWDQ0cisziMHD8CTjc1Akbmf1sOc9fg6oOeJLWR5rhQU2nPiq6qkYRZ
42MCXexQQPSsXa6SROLHKIq2/91YPoXp1jsbiHPsoA/sL6/rqL5jTsRq1ol//Xu7/OLeN0iKwQkA
S/mcyIplqiksSDH3/qufJ7/sQpwgVEeOrNy0DDM/ga4i/FQRzG40lRoRcRX3oDqo3+HYOrinePfH
4x8g8x26ggEpRBP3xMTsCHKPnbc5PeLRuDA3RHa8mYIOSc00jytX93mvXFFYgL6A/h6ETwoGlNJ7
f7/31J8sFg55nPjiGQV0yxKpgkQWFNwGRbNpQi0+ht8J3xqSzoybpJskDRuKg+aOjKZBztOAcqyM
0KGY/rUvDVJNrVZp/tHvLLzwjhRhBVdZSJ7Hv9+VYBXVmqpotgh139oTFz7PogE7pjvYmdazSsmO
fG0EWpFfJQocx1mvR33GLSs2uyIAWdbZ4nedz3UYbjbrmrHl1JLmvfNV30tX8sE76K4hUEYu5zFV
P5Dl6eMY+efLY+jSyf/RwVozyqGIO1FYzsDx8/yFpDTa1Ne8s2w7VW5v8D1Epy8xIEtrrc1TTL+J
FPRIhpTbu96gzovklAMiqAaW45Rn/rnftlG3yRxIYgjNcZg/saV4Cc1jF5G1dMDZJWyTKFdInZRt
8fhE7mNBKr7BP16L7AeDjIj7/G2x3gz8K/MnCjUhG6QEPKjKDuknctf1Vq/1XU1jrPPdgk8x+wRm
0f52xdo7wQc9f7hkmiGWytSXoec1oOFDuWYfIzhSoHqFifDltCDD6yKopKTcJ+AXx6/fnGjU9JfT
9vkcuqQehBTQ3qMvzOqUPKK2L4EVyzdD3ORUbmgAT0HnI3BOwZXs5JQ57S24H4HTudlK9Qwdwclq
qohEuZQM549txV8vjJAR8jz6MfQVWvAU5RTLsXQNUkOL4DxhHU6KjpHy0lN3nsAcTrsVeADHuzLo
PmVr5v05nENPMg+gDaxznP54xQNz6qVFh0Wl2wzJupy5qDXZ8bSACCisOnxujQUTkbn3edbo8j25
O9Tu+HOHazh5JUYKg+6t6NB0r6KjH9HtzOjj7hDhnl1gSNsK9b9voZxryWs72PlttN2ppRfXYFY+
q0xsw6OhPckEi/keMn7LDhRVKY59xdeb/Tc9+HmIKDJZTUd8CFzdgAqHi9LwywDPzgXEaz2iJaiV
iXWfveCGNHocef6mEZJZw+8A013Ku6HwMlVlco7rtbZQJVfW2pYmuL2qrFoDNBT42fy0mT7Z1Zwk
0G2dkZdr2RgLDdEcflwr77Nts/HrLPyNFYRT7MgebZ8cz7/GO9Syz+ePRN1Ht6imKxxnMRidagNs
rcLX3uCKh5zmXjCe7TCwKI/cE7sUo0lRDyMI2mxyCGcZrVQXa8pVXZ4x8j0o474s25E0ITfAiQP1
ER7mGNtmxVvE1vK+ygcCAVwNlWAja9KBw8Zjm7hcqUydrWlNDcVFQA2k3jR+j9mwlqbCk6GBoKYL
YNbFxqLmpb+9LwmmQhtXrWS/6KtoRFCUGIjBmhFFgmZW65lzoHyLrt7/NNbkEHQYjHghjNgPF+n+
viRbDcj9YkYYhyRwutnlslgIdou8nmykW9dwqvvQPMT3O6QPZsyY8tGX+QaS9V9WtioR01qwThE0
/vbyA0X61zan4gvxj7TBcODOneMvjJlWTw5R7y+Wwfq0NXKqXP6MFaJi3MdAJQIyC1QT8sP24kUs
voeff0w7CcIv6RijGYZo9WZfJCnmlYXr1ex/EbnYJQB41RTKbEx3Q5NLr/bHcTWVm/8YcyI0hBqk
o5UTUJDVjhPc/E1XQYl5hvh1qjJ5sjuXKTXVAVgDknw+0bMh746u9wLIIsXbEdJ5ZWw4OEDiiUBO
j+N5GEpfD/wE3MCIjNnORwBWelB+1IDRm9BYIlqmDnDFNfCnuz2QADE/nz2NYBLB6BqRJJ5sQllc
fepHIFNVPdrCVBJYkfdDzBEMchozxo9yE1iMXfT4k4bYnlieFpBSV6EkZisytjBy4d2aVROy+Wx7
zrqqoBqf475G3W7pDhPWr44ZAgNc2nxNJzJOKrYBbiGqN71Nst5gXl/ZEgXs7Uee4pRno8pxByrX
GCv8cqW+N2B6l8G4UWDV5MM2HcH1raF1EUUUX/b9bquLkpmq7E2TiuQGnlZgnZEqcbzhIKc/g6uG
6ujHjXtVRYB2qO1t+0Xt5+4/DsLFvQIZxS17wJfQrp83QmOZyJtSFhuGFIe9qcJIebwwZJB/C/wx
I6CBawv5FWR76dzqcAc78j7xqxpDylacWcvQai2xjRcfAF4KU4AlTXWyPP3ydHs8R/Bey8jF0KzT
D1x65Mhkp21huoXJzb9HwuF40vYnB/ToiJ6VUVKUEVYsbBtAFfi00Ib484oE1mK1jrHvSJcADsVV
SgtQ8b8XZfHpxTpP3hfnOmz4fhk5wskyeGEDXZI/tuEmGSzV+ZXUowa9kpRe1tebREXytM168FOo
EgGaz6YXbV85VtPu6Mb7YVMDoEFdaUMfUX4vz40E1R2Gnk5leMbG9vog5gVymr+hYqIgwdzYsptU
7OrLUpzXOSIgwfTN7SqYDwXKYXZqnvPtYkTYtGqP97hylh0nCX5/2qACa0X5zb4QJI8ijYNRKNrN
BN8CvzKK89o+8lT9WCYVDcAAiFDjyqd5t5uFFGDZay33kfDiz6NHsx66Z+KWOk68dhfhLBubOhh5
fHtLJpPL3hf8ebiA9JVtdta+ZwSdOWEfDKocBSXYBBrRYiuOTEjP7lQKd8oVyMZQ3wM+MwQjTl++
SdjYUJgFHiEZuQ6mTDfqQe2K5tI8oCOtA9kXM54XQ3gyWNRqJPQ7e9owJ3HbVVwHTwP04ZytysrV
vA5JLoOHXHBTKuxR0KOgPGxZ1wFshiL56JdJ8mm7muBudrXcJM59Lzg0oc2Ns0tygfC/22QNUwis
cl77cf7lii7CMmpJ/c6I2ZoRs8u4sKRzsbXQbqopUjH55Hksto2A/S38i4Iewj5lZoqoCotn29sN
jDYwQPX40qYF6qIBkyK/DhQ9EANGamknKrf5EyhZJSMtCS4tNpx9dyIXp9xDJDL9vYROQXQQEb8t
sH4mvd0I3/y9w+hfdMGDFgB8xgxghgTKe+8a/sEIeMYR/9LI6zFUmvoUBb9T7c0PlagGAlsm4G0c
a1+n+ukKYqeJ47vujTjNIopAVEdLUjvJ8Ticj7MrreZ4vHCsvSSvaNioxXl7sUQhoA6zOJDhrhwl
StqHoS+8xbUy5yYgaYtulvrfTgQWmkEz5VzchVhmKkiJj28/kYXhZaaiWQfy4N6DRDJl5D2AVqqR
Mm+2pDISwY2cJsYCt2rpqhXeE0GqKAHmLrxcJrxe1iSI7KQLeeJjlua5tEVMjEEVdTx6kRAEnDBO
JlmTG0ypzSZN+WoYDuElddFkBgqEBQiaZAwQdzozbBnjimQcg7Pqi+7RbxbRKCop+PVo+Sgh5CMh
X4jnw0e/JfMpo2XRN95U4o6deYRoYw7aFczjNhVmPltboJ3OW0DaDLSd8VugS2lTaet9KM86GPvt
YsiMgGBybFX2sbyPtwzzMgpikpp12qIoN2JfJSVl90Wno2HW6kXgzE2m400R6wMMP5h9ZkF9dwXx
bFURzARBz6m0velBZG6eb64S3pg6OlXWx36fOHV3GRfzHy/FXqhHsjaw4k2QuAAXotZUXHNsChOl
E3DMxSU8mxd2n/v67la9cq94zQiML9IfppDiQ8yi3Zab4Uv85kCiY3p5chfwPbbs9goC0Y5+GM+3
OgW6kVZhq9dHFLK/91+ke6iH8OhfV5MR/YaRHLd5EPYW1GXgGAsAyvQJzEMAitMp28V15uXcO1V7
E8E0p7/KpYNU/RYev7Fo0ttL7H7zNWPUpoIAE1HRAasfNFX45//xsI8vFCjupcypxAJugRkmtB4i
+hLkcFNCEKIo6CDzncaoEMzqjJd7usnHwyFZbWIbxuz9k1ZkcDXo9Qr46gwkPdbCO5YtlIgYiYPC
Uldy/QZa/Z55gE/rbJf+mG5moEeuVWg4YUJysH1ecuwqk7yDcHR8sG9MsvhhFWmmZZqHnExSq1J6
KPxgWdcMe7WbYjTSkC51i5+LMj0RCxMFp1H7xg9pITG3m6J5MCR8s5nmnEhwL9BKn55gK7L3yh2K
d34STmPzq8otCz/GyPXQk6DHdmVkziLRDxHCswT3pM7ED7qaQQYlUr/LxdZo+WDK5LW+9gHl/1YE
9G/uQpXz6gnv3p6TxUrMIrL45BfEAUVJNIp/d9kBnjyEq2G/ETaqPmT4gIUiFYJxNIbAjQN8oMPh
xzm+ShkAuYMp9cObU6NfXC83kvQR9YcY55fls9f4ocacax/niYCZYPkvkzTVm36g0kOROBu8Cmb/
TqNPUVSvkUVu8KZN4EhhAwN5a6lvZcdCKDzWDSUaeJhQsQw/qSLn1vc6eZPnzlq8ZlS9fBQ0wjrS
5RZPB+qD0OGeN3WatWgXMpLmxwP8BFBAHu1U0A1vuPDe5m8iR6FSAZbarqEKF5F+frZyV9/6M64M
a9XhN+a1FcmlyBTvCJqpFkUCsmxV6Gffl9DXyKDhLd4a+UK+7lr1XZKKchXbu9tqpVu6NoezRgAO
KfERqAYM7ytxnpVdfk8NkER4RkC+qqugJtqaHFP2o7lSbtIbqrOgZL6YnSTaAR8E5j5fJ5IkMKlt
jpz5mYfrGRa6LAWGQdiYMIQJJnXCTzbSTVeSniGP5AMMObfNzaCqOgGgCkFBdvHuJR1ztd5svdO5
fksMTA3/ecRFSd1kfjjp+upyU4j/8vrps4b3VhwfzOE12eFx361rEEmO+ecyeGMFPbdcYWcSvL47
EVc+Ui4/m4NelzO9b3j08CSfBnSauewLZm8HqYzbXOGez3Yf/mr+tYRi0vwzXNX/GMbXgCHo5fDq
rSJ6ubbmwzyg/ymQqpulYoy67FAw4PDTKoEHLtCaS8DriJQmXLduJ4o35YrlM3qRWf78CpJ4pq1n
3Qm0KdEUJuqq8RyIku9w9LpCvZo5tC7l7TmRTB6D7bauII7CvuwdjjWHDQppwv4pZVXWvrjKpCoA
OteDzuUysRu018ptQhmzkyZw8MevZaaWrthNh4oQwnXCP6ajf6oxIDSE3dez1q0FWkj/7HhYBxBw
bdg5HNqoyU3O4asfz21IISVe61s0GtMQGLxMzYATtvcNk+drpYb6dP6efZqTlDvutIqVNVgG6HE6
bO6gQqE1PkcNivOHxM+aZ5Ph1ABF79m/ItSwCMX1nybrJxiNU3AEF67PYSFXLPi8tMjOMemEV+Rx
9Y8kh1VEjkr3SkykBuMxLuXppGwg0gc7AYyIdTfM/fcPukMP/eRKQ7qUHmUjURSKgJX/qw/8dji4
kv9wyHiTUlBFYTGGyvLLRm1VcRPInHGs71Iv2fHoB5b30MUC+jlJ+1/PMDQeL0c8F3Il4iHi033t
Y1hYdMA4z1Rlci0L9kuYmAJeD2hwCA1g+ptr1BSrNnvv1wFtZ8nG2cQqOJU72EqSfBwnb7tJYrjo
QX7vs40zx/Ge/zFw8AjySwafUfaf7l5b81fzK86785mUvNb3sK9p5zZx62Impkr5YylXgfa6reXr
iYv0vobnm+pcr0ETtLb13ilhCni+Mfv1OHkaGNnNsJ6lOQKTiZK8qr33cNZMhIvRa9kpRiNrngxs
j2oXI1vy+sQGsmendTyEhs27pqBxhc7w99HxkZP4RooL+qFjsMjYc9Io5uQlx0QjoUCDovEAagAh
XWb6Zu35Fs5jfv94pNLLDwRyazoMY+o3zhgH/PCsIviezeYbxa5psQcWAtzJ24oyHNX7qAUNt8gA
2uFxcicVsHNilc0OH/eZ6dEdNQiQPCPJMf1af2Ysp0TOyzleDhiDHHzfGlEb7LVnK0HpBNBliu9s
HZpD1tKLAkQC9+O25olW0MXmxmBP4xwNEyiXh4QWlOAAjjUyAOfPvPbibqKQOEmHi7wHiYMHz01q
RISEfrXn6CEcivRXqGZIUEqopD27HeAs1Gk/o6QZMQHaLWrYE25BblSpTejrXOwibWOB+Gx0YFiz
lRD8ZYDLIhXDUvNI1+Ltpxr6tEZe0gwVpkr8s6Ii1S2+tJZ6Y6ET+pEzUaYumVMiYxPoCho/SUaq
ZbWh/h6tG9kuSwxRSxN13mokWn+MLfYtLvELwsAsegW2SX1hffMoo0gHaZ38HbVY0sXmqDjJkkE3
NSCqrQZrTpuxsNsETD4yDSvaFLP9FF2JGIsDnbjW9cNRKW+L94cynUsgWbC8aktA6cDC5LcugrhW
rp68uQ8ZM63KjdhGIAkenvdowEyyh8nv9nPAFZd1WepDuY5VAsQfGjmEbF8CHkaHSC1yDA6cZ/AM
dtN9TEvysrUHTwGxx+uhIbq5+XVo25Z1/7MwKtwkK1qRykofSlQlAkrhOzM4f3lLtquB1S82QoWM
N0M7a2rLOSrsY901N7g+4bAzSTeIOr2UcYuh2l8JtCk0si2khEuBhDvyC2jiHHQurwPNtb+XEVEi
PweU8v7y3CIDtVztNvHvwWu7H9/SJMBW41uoMGwAAaPTqphVvn3fnygIdPckEIKb4lqTVGhEkODv
5b4RJdOI0htDOerzyQ083ssT7H5PdDpEEQSSrbgngmkVjP+GcAfW8J3KRM1VBredTL+1Ck0Dd5BH
QIVrUrnK/EV6U0jDYZwMyuqlukwxcuv+m6+ksH9fBK9BTkGVqofN/EoFciwJaiGkB0wd6glbQYYv
EKDWtBVmP4y4hX9hp0B4MEIt4ADgwxN/8asGmbIyIVDBXowga5Hm2etToQeYE/F2liNLt2/sidee
azosbCbkCft4orPqWYEGAZNpLiABySkNY4bgHwNAjZrxrJdG/jUhHjdboOWxJZjli0N3UsozYpd1
vmQjhlvwYfEKizkhdDdUDIiXwDxGOJUVzv/eyFtoNp2dBxNdq80b44YuSdpdWqAIoNYGfUF0W5z8
1h8zoDaV/xahhXvsdm9YZo5NkulagikCwwg1eTKEdwOH28QZP5PjtWi+uSNvC6+ABYXPgBTp0zDE
jDmjlKH3hnb3R5nVQM3ZFNfwUDATcosTnZ8X9I9FGr0KPhpgBCkmflfNVJNMKy7aTnLL0KI0st5g
MJRj/KrC6jf+da9bgE9bzXFsCE01DSdh77YRn5sctxM3ofaoqdsIi7REMvY3uqz9EFW8YLRVKcoE
sbsBy5BfOF0rUpKB1DnPY7jwgH39Mini3P2DC2TE7w0AQ5JZJlm3h+O+EQyWr5PHG7UYtgf4vKZu
7m2P/eInl3DHJqVhU7LiM6cyuamv0zCbbHFJxvNgJSv0Irmv8YBNCINjWC66ss4gFU4hMjo1WtO0
B0jU6iQC+Z9sJgPrFDnCZCkwyAd0LCKf3JYNODcM/dxP0GppbG1K8i4F4L2alt0CVulVZBuUdZwB
mwkHsMC+tfcv3wisSGVfUnOXZJ3iFeGVmABSQ8Xu27swDxsQuvXdW2mm7IA74hSY8vVbaoIIvfvE
a08OZKr+eAVf2sulZGMlRv29C8mkiRE4fbXOKD/+ZiBy2FvxQgFDeTiKg2KYzEM+V57grUQQkXPC
dXJt+/LBHcC3N1RPjOzs9uNbKtiZ3CU0qgks658Vy65kX6zRF43+7B0XSNUyvo/wN2NdecX4cLNy
RZaA5dNhykXxwpo1X3ypON9rx/h4AeBZnRdqpaehNUOIAfAiWzVGacF3+wThTlIskOnitwQtNp2L
S8ZBAPlxugOmaxTQR6DNt1MwlVdWTqHpBJn1xntILEkREWUriraxWKW7dyC8O5epFL3f0C6XpL39
Bb6RGDUI8GpcEnFPvSwI84dnNkiF33c9i6aNKiOr+vrwpu2mkKBlvfbsHz44yYfnJFKHXDXM6Jde
jKX9mq1RaerrQE3vtvVqsf/xJgYtcYRvxiV0pRvYIghzi5HXx8S+X26i4lJfKCUs099SwH7fCU0Q
LXgBMYC31gVdYHsRLhKfUzcXo6PLxJMURFG7y4x7tW+jZlgJzMxoUyBjRcH9VwIbvCBZA4LGz6BS
PwdJyC62zhtvbzWOLJUb3+/YFcL9CS04mcdpzzvlr3PuVO7sl1c2gdNkyaZHeksDnxG3lbHgkBAq
eHJVcoBWM76jzJg+bQYzXvIecY/znViajAb+KucIGrsHGK2Dey8XoNIN2i9ONwbAKSDOpSqBq5XW
+PfiMXkyvImrceqqtUkQMo2G71sUMQlTV2978gmUXaI4Fbu+tM8aiH+HxHGUqS/uddmdIY+c7ckt
VjFKMIdb25wWnoodvsJCQyfBRi5c6PvHR1JqKtsI9MOtOzIGTYMjELekcrNek6QLgnYP2MaFuMX6
iGY6iQXRXjPnUccijhfDM5wXiaVjLbDu1fweuzR+PBKgJ7U/zRCsftybKIkY5SCTCkzeJnTuXLmV
5k1SWTE2rthIPbz+ffOqhT7Q5YeT0HzX5xa5bTxSiXyAh567vuZbtxb339mIEO6cjKoEN35soxBB
hZnLPNtVslb2hy5ZrT3JBC9tTHcsd18UVjMDBQj2Qz2Itzg62HrWN9oe+kC9fa6LZsDB8wCfmbNA
/FFp+wo/D3+DU1tn/pwxUuX9XImcEOy7jkyt5TuySqHvnoGQ2E1Hsy9sU3+fyMu52Xx3zkqHQ33P
tCVTwUffzN8YSHHas3lFrVJBgHqyXfwsomvM2DWTjVo6x9tNARDrLZikvjNQHTHnL10eOXPJFwwH
2p6KV6+isVVFy+MvAE7f/9AmtAqI0NL+MAftgXaYN+iiP8DQ206BpayblCi1pQerQdOaVRMsSF+k
Nn3zyaiJtqHmopAjyL3E5+qeLBiJPNzZ6Dtp+OME3QqFkPBoPYlF3yQ6o7OxsinVY2Cr8V8MJHRS
EFDKES6PuQornfQL1T08RNc/JZa4jCv3h3w0IpojPWtmzflqwMr7pCBcn/bwASQWymz4AF11XfCU
KfAQIYCzvbGOPuFQgLzOIAn7U375PhIrMaPvq/ula+A2ncfKz6dAR2mjFOYCTmnicFy50RWpy1HQ
lnPh4DrwViXXrQUOvDlZfLOoeoDF0gi7IjGWB5CMKihLtRQWa5m+1JVP/Ox3bPD52khvw+MNEp7l
WZqZq+7ELJXqps3+Ii0tyYTCqm5hdjxF9QiXJ3Oge1ptRxGsooHicuMPLrzybNicDvx6XB5CEbAt
IIRnXKcgwIVsO7P7DBWJB+b65//1yuERx54mUsFSBCCht3kKvmKEmiKVgtnYgBTH72mmJ5ctR9YC
coMKbj4nAOvKwjXQIJmPdFgXiZSHq7vjsvG1VZnQyapmDLTew4B5S9SnbCO0NXReRZrpR5uk6Wss
YvYUy/8mRcPxSytyBRw5H/1DkwP09PmYXuZLUcrrU0nbvj1pqwvQ+L0lPanIyMOJsqTFvQBzMLj1
6p47NQp0MCu8Ss/vNG5RdkCh1e/oYYFAIociz2HBFbezX0eVEXgXJwDGUIPZ5otOvDzsit2UccX7
TKbjjJGm5AhSKP56hHNpR66tDnQma/Pei/6twe+s83KhPXjEMIN9CsgxYb/HQIck8ZamVroy8fj3
AkQcOacmGLpoLsXnvVlF7jrIMxhaR6v0wiE1Ewj5GLvz7NQjMGCZpCJ9uNDZt0RhSomvdh+EmbY0
5J3uDLG+sGJm7Pzb6PHrc2RxGFjCsM6KGum/dtLgQO+mIzA+frcB49m1NJ6CFnYBLZDH7ah2e9E6
i0bBOuljyQ+cR7AgBXjLBTDDoJYyWB6CRkxZguSspTKaeqZbWHmS5mYFapqnVO6EpUkSJY/7KM5h
LyxR1BKzAZPNMmWc3QQfEWeN1e/TB9n7H7r9FBOTvRPjKEex2lJZdtIaMnH6ZTU9zmhO0Yl+OtQP
ahqQj7jxsCxKgw0pKEI/YbryxuWM2ZncZL8Un2RBAFsE1e/hV/PrK53HDuo6SmFJXEz15/1tlfIw
FnCEiQ4JDFNBpUG14HflxhosJ2oe++Cqp/xU/xqAlmF8RJiVPXiLcDC9HHf22uI50Gyqc/7VWoHJ
6tTaVJJ2Mu0sSHbl/UpDb95bNFQktFdZjXhS9U81FmjqHjmRLDP/jXYiJaPmpbmbVBVZmTgTwN1O
RL6eBNHRUB55GC9BKmtKuWsFzNku8v8BPJscUtvmgwMLwnkDtxEmG49DmhZ3Ocs2mIau8nAX3F3/
8r/CGdIK6YhnpOoSwrXEresRtp/Uss3NQfzcvXH/pRdfKzEuEAhXecVljFclZSE4jUJlBO9xAXuJ
eofWXCxZDJ4+Xay26ETXYqC55EM3jCEIptD0Qlk2aLtnWJ6G8SZfAj2/Lgr472sLOI81lXVVJukQ
XRUH0NbEkk02/BY9EOqi0l4Kep83FPJkB1AIs+rVz393+uXuG8hPDvBsnMmf8N5xeKOWcAmM8+Pd
tdGXKJAZJdyp8y0iXVCEN30dlyTJUdMPZFbo/MYHWlsGmVVtUc+cvzzv6F1FzgF0bfyZUy/BRVZx
xtpifqBXqGUOw3xeZ5QIxlJSf9gsM0H0Xez655cezyASX2/GmLDwCSCVTYW3MJgFDabxfHX+iduT
1uLOansfdXvRVlYc6p3v4wz9wh3MX2P22Z+CbZEnrv4E+WiOHwyMrQO3W+4pEWvI1abzp0CkAARZ
hN460uJh5dP+J6bz3eKaCprAqzgLuldVAvBV7SzLWymYOzWP9vUckgq10rfMeKuiGft4fqEZh0yv
tbJIxKAf0fylXEcW5L+cJgVmT3LJr9f1b86Xo5PMuX53sc9hSaoohrsdTppBB5wfVdrRococObsp
p+4wi9NO2Lbkztm8gF2dTVi7j+jtFDmPTadJTRT1LCWsWeWYaUvVATPSpL+j9j1zo2sNo4zq/FZE
tXLfhoLDp+zgQnL9vsyVvV7auSUAXz2dCEM5dVMzPNbm0QCSZ0pAKf2etyPqjKNGWee33utQBlLf
NI5vMI02GIU/FVoXtt5oOazwYYBhaBDs2oGIBJ6TIYr4NnQDf+M56bHV0U1hUy4v6KcJBZBknBB/
Z4VAGOVB/b80NJKg0hbN6JtJ3xqnmDdIbkOxybL3w0OLcK83Wy/UFsBrHchv5DDNQekj/1SbIDG9
BODVYLVRUnEXmwOplXJ397DXeKNke9kZ+bZgfU/sJASX+9Rto3BUiN6SJP+gN7X6KqVAaDn6fKOz
m0L6sEVmt76m7S4ebpbwvGN+oQ3ahS3oKYkRA+HSPz7YJZqe7rTIh1yGBZ6OhVXRopLLgWFX10od
Ahe0hBbNc7eWmh4082fJjGKFiBeOQpKS/WGp+GSydBdERzC5LNvCKUl6oWzubQ2ZU4pGEdb0CM4r
+zL9pkOmAJmgP8kJFjG8/jJyj9kG3PGdU/UxfiyrwXgdBrMCQ+9bcTbDBAzLrGF5ONEq5og0nIgy
KQtD52ZRXztMRY9Sb9GQ6kZRKV0CYJ03NZLPaEXZhePLHtSYE0RzYitmw8g+E590wyIbVnZuvaUv
n+XoYTTTLoqeQFp4ns8YQZY0EcvSbtKMOwricx4db66WC4HiE5Gl7iJidbZFECa30OxRPM1MRJ0c
DgZRICBjVxSCnoGjoIwoVuIZ15AxDj4/1khmnWpKp1eed1OMFUq8ZXAemz1O1Qx3lPSDmqsCQd2p
w9aV1Ip+fO3a0bcfkLd9UPouEdJvhzkA1WSNO0seWJis8oNSCLoGc0v4GOczE0xg6ceVO7oPw+qK
pfpftaGxAvUbWbHSw1Vkcr2wU6utK/ktq3NVIMvFgTArGt409h1KkopJPDhXNHnHRarZFVhfZX5R
QxvtPlyzvRvW9BnRQyjbtRmJCjR000pOdDjaSLsbfe1XQ/eEjsZjoEe+G6cPSmmBKFzXCJLOAV1P
wKswoCmeXxP4DtzE91HwUVivrvWykmaVVzD2EVIUo4sUBHPygViNmJ7B8tW5QRswWz8Ec1FTBR4J
9L1vvftCbN6EFO8+bCNq8+fjdK6BkpaiFBmijIwIkJ4cX58Yh1uhxxkCLYjDIoN3JU8QZZYDmyi3
9jFbAwciiGocWljARuWW2w4b7/Ij/gY27RYqLxbxN8mB8HASHmV1saxzYgzhKv8c95xlZQkWFO/Z
F3sKW378M9uOD+BU2pa3GbFdHc2q4J2JZC2b4LNK1R3xpv3eMgMz1EdxMEQ87dLFwR08wyVM4tSh
ckIEAxdG1K83cj4R7IDEJfK7NRL4q/o4eddApm6XbgLo9eIJ3IrNlqQSEB7L0pCTrXCCu8xJQdek
CAgVT1t4Qwv9deQhO6CPpPajcPuW+No6hHaef71dwqs54fqmCCvFJxwOuRkXIymUuiM7syuzS94b
4Z+8wqiYuuuQXc1TcvuYmYWS42h+5aaP2g3Rd09ke7zcCsdTvWQy3OfaGDlwvrUQNk8tnOY5Y0hN
pmWKpduhrl/3gSeAUraAGZ3YlK2yMtP+YvLGx9CzYVMcVPcV0/dYgULbRa+lIGarpT14MicrJijb
Ff1XSQatFEbUfkGodMN7NxyTfN6Z7LMk9PdJ4V6QSScfqDSmgha9EeCx0NF7Ca872+6aH3c5rCM3
ch4z0yo3uutWb4ASiaoTTpdpuxmDwNPe09tg2HcskU/QUuGRzvfrODelBT/a3DM0QovnXLZuLW9l
gXyi8OLzN0w93mGwISE5hmcis3rqk0DpaGlm+dCBZehYXiS/d9oe01EQ7I0BlJoDCotF9yuUossC
bKI5uj4hA3fQheM/xY6Cf3isIoi5HbqA6rUT2E2ZWqz5y6UQmaTdGrblTaR/2yn19tEK5/k5uXYd
tQY5idqKYYbIbjk6WJTqd7kWNVg9lqkju4Q88QlOInbrZ6EIXrn/1D5sFoaDX/zX9nqabJH9kt0z
Fy/YBszW4Mj/HS+QsW+hfGd10lUUOlo1rlTMp6eKElGvo+s+TF3nImJGCVN0eBqso0RexGUh3PpK
w8RN+hDQuZ+1wlJJqXiejXpkqt6Sv6uqpA1pZRY0gQcm/NXZQxxzL08p3fEvQ69BjFqlHIqnYGFb
ZOymjjgv2bzgMDieF8u7MlXG/eCn+5aRDhgQRSW5unWNhhoXsAdmAVKoEpx+1k5Ttl2o7ATqXjX3
m10am7kybV/cOsGD3wpVutLw+rQKiJXdGG6Pj8CVfUE4eGsgWJJNIezNM0OpqXS6rxb3BsTpldEK
PCMu+jcFWWiQgROfzxg4ZCqT3KAwDezIaHNM8b0gh+5z641hWeoRu4tnq9MTTymrj8KhdEWNFYBd
NCkiB7GRauxZm5WJTu2NXvLkMTfTvzwg61YEPYo04vgQPPhqGSGP/bH4jEjXsNpBNhsBoGryZ9D+
gKslZhSVu1dbNeBtPOgmm2oOBcv0Hh075SS2pE3N8la3SSSE9wWPraoFydUeh74IcwnD7krG9huX
IPx74i5YJWjMTjInIZw9fKAyN5oRW6pAKZGSLzGwFGVMX8vtvYnlVelQuSNwrVJD4z5A6iuYt7Jc
Q4eiRAiWUnV6t05HEIojOtB9HIPRxvVNFLEj4aVJClufHlzN7NCvNiwv0q1qZThWVRBk2CXpW36a
njbjNZc7WTY1S7q4bbAHjh71Pr0Nt5Rhn9RCHPG7Sb5TDy/HJS3b2YRvygFaoweiusSTHAks1hG3
VX8sADC4/Mifr3bflYGjlNQ5vnahtfD7u8LN0f4gSnhDIsl/AJbvB+lb20Qzvcnf/5119oUG3svR
gksApYzJPxQSdAAV9sqT4aWtMIrr3epS0Q6YmLYR/n/f1v0MMSgqvv8QdqK0dcjJDrPSNJKDW4Xt
cSYYSX/vmzancwkhyM0c78apGsC3ADm2v/kJY/doxq+rs8YNF+Z2Nx/F0hZw5qB3bFchki1yNAUE
csz8FwJN32kTxp29XaRIUpP9RqCz/giCgbDT7iW9bBd6ATmFod0JyxC/S37eHZYpUkmo/kqcC0aA
sDCwHrBEy9cBxg8orMbfJ/+mKdpcIGerw3panBoZkipChbtz3wdtWOmrBkiFg31CJv9mjr8mnWpi
ohkwRTD1PAGq8rLe3WZG0GD0EswJoYqT9mRhl8RV/r7B10Pv68rQ+/oyNbJYiNpOxaN7W55UQZLe
yU9WlIoflyHWEKssrr4LOMXSvrBUUgfll1seJaOjBX9g78BXjzyTuzFOxrTwAOWARrMMG2T0Pu7E
paxGFAsR6BT5ukCk5te+IInfyKIv3COh3MkFOVSgAcJA+ybLB+dCv++xWNOUslmzeZ+uoFAKfax1
Y6xM2Ps7MaSgtq/zbGLXGv6Q2iWg90HsQDw6x0nYFEP2fAZmkx/VjO/sp8UBxbQQube98HDp8cuV
lUzDKPwV3uW9fgfHju9ys/W20A2fDTVWWPzxzZ2KukkW5M14zd4qVcIZIziDBVikrojvpLIr53HG
733agvAEmkO11D4KPWgbL54Gf2v95i/oFLlQEHy5OzRiwwas4WZW14crTdUxCQPcluL9RtpLWdLS
EPlsS0E7TBzkDhw2gxpC6iU3GF9fVPyWs+zlsq6ba8lLGUGCE7KiphyNOERtKubg+aBVI7S+WPgY
le1kKyTi7NzB8Ne4Hmlud0GD82KRUFylnIwvLtlqhPb1+5pLqVi8+UtW33ws5k5+iOf0AAlEyfRX
PSyLVxl5KpFKpsDfZ1fifqHjdz1ArDXD0T/bvGhSRXGGfrCt//INL8D8UC5zkY8SMI27uGHvRH2V
iW8SdH7EiNvDjdb/GEgBwU23AqJ16uvBUi8hKrCrLroaQ0LdlOEfxlpgElgTABil+zUXMrhY/9Rb
BUhSOC3I8TA6e4+tgpxJmsqLRrC+GAm24RXP2HTK/df/ST9hIYNw1ki0LakSAPPtZLR/L2of9d3K
xzxUieCh7HcbYr5HV7mIZhMkayWnSW3mrYpkAVP9WWmersLBeOOfnB4FsxPcnTLLFaeEgDgWm5H7
2YRFPmOoyhrpkvJuDZHFZe43B+n60eoXxQGMDizMAI/JO6/s9f4eMzGOQuA9MLg3TMvLskZp37zG
zkN4iiQk61eWivIliRmZx8aoRD+pOsR91A/XybATYvbk7y6xhRG3p0AzGRVRjDyaQ7YId3xjpYch
HYfGHMg6tj0Bc9Hs/UAMkTjCRZ/SoVlbC5wi3aBSipCQQVTnFwozQa9uRHEYtSiX5zhSe96Exwf3
jXHt/ofuEM2Q5MDiy/DY4uI39GF/uAuVDSFpQ91YN25v19xh8LEBHMLtGJ56H/sBEjg5Kkqk/gZY
nXHU2VAEUraShdomgfu1xdYIrNws6KiczcKtnOACqhwlkkRsQm3sQcZx0OTr/NAqb6OOMmmQ37E3
xGvDJjsmSuzi5d8fCwFQ/rL8Ya8igzFd4/13VPvLwuVLqIPromcFOvforMHp79dJN5c4/gfnOomY
x3i4xNDffLQWTtnXA5QqE3iwMKaM/jllnGzbaWL4UpYInKYsSQVa1JvDfAIW0OChPlt+8m8PKvj7
eb1n4JzWV5mVQBZWBtN/of79EcgQ2LYKXGwdjcIoVFjuIrEY3081yB/baJJnuO5Qjn1ZxwB31NVH
bb7sq09OsmumAe740WekL9ROZQDsKjQFF6BqYpd4ihDHeLhcNBs40VqCKzYBDiJDTVzovobCbEwT
IPgMl7bTBvN4mx4FJIrztky8BcyEd68l33EQNEd7FYYAQ9R9TtDjV0POR2j/vB36eTcS2pcjrUbK
xqKXMxUfZAxqs7E5/m8Id3mLw9B8IpjA7KssR5HIiQq2dUqM1nPd8kSQa0UQw++92l7LV5Z9i9vu
qsOmBA1kTpsm3n0E2Ui3YfzDvE5mXVsAYGqSsRdQzIwM8lTsbb4IGtVKIMx8DmOVqeTW55cr7374
N5rzJFOKwShEvg5Xlbl4WqUbzMVhsyTxT5PEjEr5lchxwFLeCkcGDt/Ua9yJ4N9SghYCdc+qEgYy
OX5T7TIaHh0Jw42DYkKjl/CNh5n3iiywLVk0uu4C9f7Opst1OTP6hwHi55LPhLjsLHkOP1a+2BjQ
e7fHilOheHpLpTUNz7aWRkNCyXwQ7BLFmpMIb9NV6ccUTFlYiI8rrHqMX9bnmgfGY0OERCLNrYvk
P6wjvXYj+/eC9QszAorOMRc+GTKvF1klO16gNxotYRSvw4ErPL4sBA29T6Bn5okB3+Hr8Nlauepu
OBIMlrpuVtrE/zGpAc7xU4AQloqVz75KlghRJV4zxGnzVLFWOoBVPXRhZgtC7LJyMSoRECULrmM2
kPgNbnhI9Rw7gQAifgJwNFIkqz2Fti409OJhA82qW8FgjbV0E/gPaf889hLeB4w146wvYNx8DDXl
WEZAOdVu0f0MRrN7Qnykb++1YH6Ne+cDtTSGGlI8WFuJcyZACebkI+YppRIvg3uLIB1ugpv8dEkT
TEIXjgRvhTiFnhXnI11CQoPHsF/OuFj7Hu2YJoLAv2bGssXk68V7WyFRAHUbaZVN0US393HSgrn6
20v/az8cgDChFOsL6v8bH8/qr1TbdS5xt6Yf0vSAqgSVH85SgFhG/hzVdpDCUKzSK5/PROuoXSNd
TsJKGf2nL6KaQybyMr86M7heKpvTvJFEduRFy2rxQ2STNPGxttM1patiNg7wScuMzKpbf4tnkz3k
eXwzUyaXj8T3w7HwA6utT3YTh8exg5Xd/sVzFGDvBHG0mls6rFhHVlkCT2mvOOQuMuOtv3zv4cGi
MFA8MD2tDLp2kvlS9ZMTdkHgytZoYbWdQlh8u+18UTkhIIsGL9vNrvA4NjkE+Pvqtx0WmCpt9O5g
ZkQ2tV13n6DWg1gtTUEyy6BVGk2s4iMXUCng1jRKslbLBeIDRwAImETrPwqvOIjqgHjJw4XAjus3
v7Rg4gGZUeomAJw4ICe/lheHUiLA9xbXf6yA9pRxhOGJV4wBpe/n3H/26An5ljru3L8auLvcT8DQ
f/5/HSfwYrPGehM1BBKEje9SuJKb9SGGrp1Zywad1BDO+qyFBlWyJb85fOpieM5lTv5m84Kji88e
bz0ix/4eCbf/rAkoZKO/OguW8rvki/qOeXar4FFFiqOvIfsCYs5hIytMvHn0F+ZFiuEj/NFiBHyX
E3pEB7zd9bXFzH1CMG0/E77dWtystj3Vsnyo7LmGnQ+Kk/Rleuzqg/CZqd8hI+69/dSqoSeVGJtJ
5q12rRR31dnxxupWLgwl/6Yn7D4GPbMzbTQh9kmFfatqDopcesMBtNYoY6ZoYl4LjCuqJQ2E9jOQ
3yXYd6g4y2sJwFYt3r1pKabZJbjYAJGp6tqLSDTkJDNAlEf9qijDd5lSOxSZYjeLieXgCGP2W1zY
JLsyoR+rUhoRbYGz1E4BOtir5LH+H20SYxPJzk8nIRHDwqVe6gR8AS17DXTNxdMqeXKkt7s3cirL
Dcvd0J6MOE7M/fbvYLYlwlns0yhE1LeAd9KejiQG1w1mN1ThRW0LStAO/fotcnZgcKXVtGgiTeu2
U9CWoymfAFQf6LuOa/eIe6VMgxGR8xudoBSdi8n5ECyTIjFZKmSICCtF0zbTEiYMUKHkZH1CQSaE
KxfsFL2jS1c397i2fN5tkqddhpb7KxyYuD38qXW7TuVMInYUdC1LlL6D+I3ImLO3YcKpG9fbkozS
IJ9HEAR11yaCX9ZyDYhUdGirsZu8I67TJkONhMjdEuYqNKFZvLHHHJe8pKqEhdWh0qj/ykd/dqY4
wC6ToA7hbLh/0QLH76Et2HglnD7oExOQcIkUbE6yenvD8qRgqjTlmXsnCl9Os9hqzL0mDORO8xbl
cQkvSVIXT4BPXAdYKZ0t5rwRm+Lpgc9ma34FTFOg6Zw4/iSUkIeC/kX6hmK7+5agFBLcJwAcuKPg
mSuRti7+wn9RWnq2CmxgpsqCYAgF9gaB59dhlOgjAI8fofa5amGomTUnXKJN3+dek2D++GZFujwJ
dQc1WNOuNiXKR424eU6JrsAATGT2673QohaK4yGu64qR+7TgVmxt6WpNoZAO4VWul9LSQtC0VBBT
vNDZEYXaLX2ks+07y+tCkaWStDSBPbdTtT0NJbSGvMLFtgVbg5WlDBxmbao668fIGCsV1XRqFdMy
ENf2kbTkFfl+JV3q1zQ19aiNXcRXJgezB2bau0Su9ZuGS8tkmRP6wOdZ6Lv8HxFumPQqSyK7QFx9
LDSnkThuNW2ueCOggq7CQXn/1SQCdKIPiKv6XKbCrZ94wOedCak/6cY6L7he2n3OTS2ecj0yBIgW
QvNgkHgsKXCCG6dqKax1D0G93lsxvmEZOXnGOfLKSQ05DX78rgXN2dj7DJymXtaDcZN8tWZ6RWlx
0QsM6a5OK2kjSwhSnlVDf5m/w4W/lLlLlLbvGJ8WK5m22NULlsEU55JQCnlD0jdK4NabrRVQOdaj
ZczHYj2vcPajumYA3Dx/IPh1zBjAu4C1pBaJbZRVFhjq24zMhhltVkQRiYFUvao1qjdJGEM0tETM
Qaql+OvzBvXu1cl01nmKzRTSSi7a5//X1I4puXksraNnMfio5T2IfF5xYZTuRdKR+DHxFmfwJQmf
PoH86ZW6QEY/glHNH7wULPHk3tNL367M46Re2X0tw9WjmQXpaVmoOGck522CtasyI4M5IMonPExj
wQKrKEKa8mRfcOXSpf8YYhFa0ZuX/b7Lvowj5NxICLKHZ9HALiDcH5JfD+FS3ldFybqDJm7wqqll
WOZt6vzwC0bDIFEM7W3LhxX4t8hqrrlxUr5POMIAQA2rdnlyHmlMkNorQ2s40uO9tTQeIWrGfZz+
mr6GrS/Y1+zZAeAA1MOAMHsbCD3iZ5GQ5sglfF3HoO/kQ7YmglCuehVCQMYn64D71MBplouEm8jX
wiXccAkMJM8OgA3wnQlEMLGPrxt/1edErz060g/yrLmjT9gcg7wlxSJY/E1e4DY85nFj3COG7tGj
1sZELoCSYUToHYNubXM2T5dZaLoCoe8JaFPIJ5KCFQt+OjGPfrwK035onTFIQ7jNY8Dmv7Be7NtB
pJ5Ef0VjtiLjM424jD2rexeX01RjrxhvbLd6OxzcnggrzLdoDzajegyiO29oINmZpe2loWt08+Qp
2J9fuVlQUeNW0xjnKP/YtNNPQmD8UETtXF/bz1tDDznUUvC2+Gd6wGsesCyLgzEeyRIs3S56DK0T
sanyQP/Y1m9PcTkbSsv5oGLQ+76kW5KRptWezMsIXffPLQwj/9rZ7NoBxoJuZJec8t+xS43YcxyQ
6nOCFL+3/XtKTE3WSdh+yZHZU4UcpnIlN8SFI0klx/2BIeQJiIjyncReqgTqY7H5JS3cZB+c+32F
W90616vWGjPyooFNy9I4vEA+4Jc390YyB7HqLRhbfXdaE1rsrJEkR3jIUssQRIQj483mhQdnftVd
XNK1+twr9zINxFPQZALRULCzMYFGZjJlMjPCly9Sy3YHcLu4aQzb7amubp2SMLqbWOCd5D9RuvoU
PLkAVF8uNeF1i8Kd/ZRNv4mbY69H30EbQ0H2k6kBBsdlgL1UxreYLgOHqGWHKKFkVYwV8BYqfiG3
8oPnGGVI6JD8a0Q7vnGAC7jcUQGLf7hwCju+rx3EAG8C8paR7/GYtSo3xXXPUEdwzHkGnR0OLiAj
u5HBcXvb7a1iCQrgAmHZoKnjD5EC69wy4Cc9bSBcbqyg85Lorli5pPTvsuNyIzsq0E6M6BWibuBm
ae2lik51U4yG89XbizMbyEULGhuWow7Q7I3h2IIIQI12pjXlbptXohBgP0335teHmiqSL+xov4hG
dID7dJ+420HzTitSzZjBY29NPfR2oR2oB+IMk39Fwn+J+QVLJR5xqdycrXPV4tzWemU3fgI17wAl
yleMBAQaBYyPBCnIBbVSQcaKN4NaJ+1AImCEjMIfJ7wKe1ZWTrnO05FuC3wU6GuAb0wpbOxmm1bt
r57I5yhuG+e0RP8O2z2WJDvteeJeflOkxd569NkV32dH3F/fsLb4qokEgdXq8d0KqsZLbq/Wg5ox
T061chtG1SnC3K56esyK0XP0q8l2YXik3fYn4u+N3QeHqcXS2NIR8398OhXuKs/XPTpG51fY+5ME
NFcOTPGiUyAMLRs5wu/FSn5tBKAVNyPKJSVHgcl12hOsXZo1t9ERM3EoxsBqAA4SIDsWmDsaI52I
swTuz+3U3+FXrLIqED7R2U7R5SautZCzt9IIwCH1YeH9m/0ZM3meo4AQGk4zuY+zABYOOA3FI0+q
rRESdohthaNyOUMbrK1C09lfqqpCxTL3GPOuZJ8qvdzK4vfWFlI3u7kmcIyfIFUJhWgh0XymbLa2
1ozY387sT7b6KQWzX4nLQQ6DtDOML0LTtFiVtNQ0iim2X5K2pimc2ysTyN7yx7XJeqm263C9nw5X
SQ9U+GTESxhqjzRTI5EB8IpDFl6D1ubsybuAYIOcUalawQApi6rSX7NCrIGn6hNMSBwbEhAsibm9
Cq5Mooxq3BpbG1S9qGNNKFoo98Dbqm1Hrn8hCIjrkGEy4XUL05YO73AKUKxQ42qu+WrObkQpRTVF
ufcxeDCzyb630zY6rcyDCR1Q0rN6YTMM/Q1CLtu766fs37oOHDEG311vWJx1N1E/2ptuh3wBjjCn
XBPWA23pUweWN1NFeplmsGD/34nyvD36Imhm5FxTukv3JSid2N6rjCNDm7H6caAt3LxAIuaf6Xwl
h+cjLK+7lzCO48ful4j2YW1xsaBarUmpiVkc8E8l0OE4Q+cTykuRio+NSlxtDxdvxxb8gOzpXYPx
A0Dx7qqPcgKi+/iy323ZT2PAN7VIXDaREPeqI0h4shDyA928T7jOknC4iV8FzHcHFlSksGyPNnym
yUB3lVW3vqIXh6c1rdSgpph9tI0Kkfii4Q4XgvE7O2y5R8AvZ6zYtGn+csZ/yve0wjTwgUKaN2Wk
LftQhjI6NOUJHN2Gd16ByJlbkwNcyM4MEPvj1Xz2Xqc7IydPAltKsvjg+3rvl7fUAyJnErwY9eyS
kvUmnny+G4og4DOVrnQo17UHSf6milrUDd9GPLOx4TBtQh/s/xJ0L7AVXDk2BHAf//fVzSKmjLDT
pV4calZNA4coeZ6M+MSeECpzyaR9PMqOtsSoMmoIg0MBQmCtS+k62wbA74aVpy+J8esm4bFps6Pp
0fk7Pyu1168icLO6ELBDyabHj92lhy9QG+G27btowfy6995ystXFadSS3Rk7nFyOKBHHKr8DLSXO
c2b+kFO8rhmh876EO5D42LE+9BZhfHBBwmHNbAGOQvuOz2sFun0C7Wnc0vGAJKqW4GceGSUpywOj
TpbdVeo45hsTyRIWcDjDlxMLM8QIvJ53fvyPNvLB8D3eoFAhyWRMtNjXmBZf+ua7xF/AfmN1Q1oR
xzRRJ1rf/1aOvzLj0wBBETHQzdCdUuxK8DvOnWnYTwjbhdfegoChMi3194UxzVsnEcc857Jzb7jp
veIw7by5GGeg7+7K9UeKVmb2GX5AF8Nr4YZk4d2g5YzlRub4ehzrsGsuIZcJIHvTuHUTjNwFwUkr
RhHFLSOr9EDIkmsczvP9Tb7c1plY4dmBQkChR/cMQ9vHLUy6i82Citb+yNIXlkYfuPSLZcC530rC
/BHxsJs5ReMbieNMEJ6+N5LX90y85735bIDcMlFu8bbWnQ8mcxBrwTZeV7LZqOIs8PtqRYh1I+6/
WM+GfFte6UDNV0Ct8xtHCs29Azxd2tFlbow5XRYAq/ctE+N0BAXWk87uiXa8t94K/VjZOIqBTPXZ
PJP7lh2R4phPtDC3J9bgRImvF+tlelDWhQZvH4F9nkeze2h7CEKQSzi+6bO2seqRfk0bvp81UoSi
HqWBG85gGRofNry06ynBcvk5wbZ+TYsygxcqxHLjPRpOy/0TzgLXTRBKO62izJTiPkhrma2kjQTW
zH9CE38JP9WEv/cvG3ZT+jrboq/TFQibOVNZsbc6QgAHTJqRQ92o18bLi+1pDcfu7ZI1XqpJSWJ0
mS8M4NlIAF85DrKKxYH3Zeybajc7JlE/BPBFLcPLcQb/LchkEks6qNqNZ+b7CA/+YvnT3CYFkcnl
XzZzN/Ts9c9b3cBaueTh/V0OmCV95VjXHP+D+oe58N8pPfBHTigwyNFL5W1bQu+Tj9GYnPI1rRJ1
/0OFI8DS9o96p51qQ6YqkA4uoHw2pJYUvkIrmp0X18XKJTYNT0aQDLpVYM6NX0v7ui9NPQTbAA3C
+MD9Gd2odz0r+r617z9JeYGEEdKzbwcMxiakXS+5i72HI5D6ag8oAYROH5uL44ykj75U7Sfwe437
8gDN+GpeIz2Ik3XCwyEgIzfHgxY8C2mUuRNvjtEiKuQwySE8sfm1sNC3mALUlE6nrvQJ776Y3AuQ
bbY9W7CKdhZXnDqGueY3R9fNpBdr1jWEWqq6eYbBodVtOz2viKyDzgKjAheeCZJDhg2gSKiFXq5H
NyQ2e8JRJLxFDiIIR8vADo2nc6v7JceqqSiIIs0Me5Gfq3++Iv1NR07r/z9FXdKphfPP0vrVkukW
H+QWtRNRVZXZueQj7Y/jBteTwYuCf5IP2c6aU1FRmKefotd+c89htlowSYgEtFOIw8rAk28MwB9y
mLDCtEJ0Wrbv9A2EYaM4/jjP5GZ4RQGYqoo7DZQ7DhN2Kt5BHgNmkOOVbYsS1GlV+9Ehvffa0HhK
tXxuazZ2oWjn5SPt/NKx1AxN9LQnQKZAuaGIjibiUyXxJgrfKTg8gI30lxJwq8aLypQbRDw+8Uf4
KMcCpsfw7qdR086IhsN4WA/mMX7jJo7Epg0FszPaUPmoOFbSyesFu9M90/Up1mP2IYCw/gIdq7J6
3bNWTxV02rw5p4xnyYUC/t49J5RCXvNy1WakbtMZxx5aO1gQzrlkHDRBpvBA6UyrZCjO9npkQ0V7
RXJXUjPs1UJghYrOCmq8JSxekUs2N+e+aIAQjV4YzLOGiFcPoXJCQJEAF2eDk1hFGxrdmp13ziEc
mkUkYavF9eNy4Aw5DH0j5p4KVZBZXihh6+0tfXfp0Y/mMSqEljWbjc8GRtmD7GEiSUh61bo26TK3
wY3vxap/ysNsP1tyY/3xTv/J00xYPDsbFGXwrCDYIRjEHSctjkZMmrBw/TmkncCxXg0LP7SEooAj
k1PuEaf3VooXjHe+ThET1SxanR/VdDADPougTgKMBIzbwkaGUa5ENxsKq9OGwFloqSuchuaiZk+G
8dItytVXNoc/sKI1DbsmXQQ2oAnlzQQejSw/wXXZEqJyhRxMacdz/KeUEz1zjpwjDJSH7IKrPoTD
qBp4TTmQ5QIitrMSv6kaFlFGX2QsnNi6dQAy1YPJdxiLZacemu1PdYWwDkRZqFCMjzvv2mt6lsvp
FbhUuZnk7eNar36VKyaD4TOL4vU/lF6WEYXqESvH9UNu+PKlGyXxUZ9JcLDZznDDH7PLNuOlyFPW
sGElxeXFgGwB2lYtIbSJ7nJWdENMwzwI4yFG6lNoApHe9DjugJum3gOqGitm7N9K/KHaPYEL7aPP
SaDwytoNb7Pi/wRNoYuygxrnHj/KjxWVC1YSZVRdIoUEs35HK8NaekePXJeFX1xZA9+W3Xgdm7py
AFjTlj3Md4LXn1mf8CEBtaBmKwU1SxHujglmmthxLj453oKU554iA/UJ0x1dFxcyVF8OxM/1TN9Y
vS3+OHmZ6ys0NzxnJgny5xvJEt1sxhrGNc9jVSD+snZykOJ9KH711XMzXlJGwo6rInD16zSov/uD
vtalmtb9i9RvWn2+9kI9CqL7FhW67A7mAgPD4lDZuEkRyUIQs5KC4UAyRgcvhk75AfoYLGQsmOL/
8RewQ4mbCGAmjD4E/SD9v9O4xsTSUBfQN1C+ebRY6GwJ9ksnI/UDvK6tcVweLzFz2naknuQx1p8h
w4l+jFvSw91IKcWi2/5WzeB+11FyDqARNyYH8YJef2+spiHQ1sF4bZJOuMgoUmmGPtY4KlZrMzt2
j2WDUYVvnGsqkRzhAfWAB29hEz4Anqiz6SqAdS8EhMv8mBRM06FQo/RGKfSc8l+NBkH6i2ULucFy
vZsazGqwlJkq67EbxrF+7Yui0Ld4xCp1NMC8n4gAy8HJxM+a+NXkpZuowwB5fSengvERte32CEj3
nAUzxDHQwZZUZfHmf6FNeae4kJhDZZAjMzRBv/30A1ZgXWlGoSHuIEwYJqZfEaL3cbuKSClWqnaL
MyJ5e25TOAsixWhio1CZDC3BBJ/wUgG8j70FggBZ0m8VRZEjH3aiAmN7ePyxbTAWebCQVvM7mbuc
20vAUU4zLVWz5N3WExjEPojkIPjG9jPFBQY548zTEd4JL07A6Ya5pwftpn1P/nNZYhifvz4yuHQV
wb2IMBEavzAb813V0GHXDtmY3loYVK47DVcC9HCXDuGsLsSqpvzO3vuEZ/LN5YmGXPPfQEMYOn+P
SkxQd5vKJjcy9Zlh2OdT1g0zFbLH/oVo7mdHm8Mo/pVK5DSv84bfmMC4MoVPZX8nes1ks/KG+ta0
PQIOID+EInjqOkuNS471tc4Shmqv5E5a3pCOEOTMm+3Go1ynVUsNnsVXW/c8K7ISrEiSXmhrXuQ4
P8zRQIZ2fvL1ZuZJiuCiqhM5oCO6+zKJ4vvaefRwgSzQYw7CGmSvS8UaljgqX//P2Ez1wUk+yRYx
81jPm7hYPaUXEvgb+3hh+KMx/YYNIuSgY/PJNkXcS/xdK9Suarzx+5TMSWaDILLPIQkuhQpjU3Bt
PkjC3Ki2W+NnPSSMt0oHE1OSDjDu1971W69msfoR+L6OZQX35ESPHZSMU0tH4tmZswcHSZEUnU/v
ctXoDexH57nE+arwInagtt0WGT3wJ2fugyIRfx3chWXx81ndXO0zQacYyKS8ePq8OWr/BsaZflP4
LzzTm2fG2g/pdiHFtNLTKmPq0QoNBQ7U8R6w+/QQjFdCryhp7BuUGJSXc/Jy6Pdx5H9LfRge5paW
W+nXodGT9GMgzYxDEub/fW5yllLHkhXzCf52JPQ5bPNCGbky6Izn9DW46AyPfA7It8oXLcQoX+A2
g8u8HaN25aoWYYXBcg+IWd+tAuYUCfgTpCHYvJYiYNn8jEStR0RvHxIs9pvqnB44LMZg8A2xxqln
1/GdbUou3GxcAgxbQfHnaKYwpzyhBuo7TKrsknZ0OctySDTufUFumHfX9dCsBIJoMVlPpLrsv+M5
uLjw5X+S76uv8ofzWJkV/fzowGUosnFth9S3TT8rfl5bmQzy/fDyNAc2ttIF+dnRJlNgUqPBP5I6
0gTOBawpM1hH33qxkULlZPBjWuZTVQ2fcRjeGlEt8f7I4TS+KGgUWEmSGxgnDTomycnZGzICJMNv
ytEAUgkRLnbzVGnWXcel0SAhK55zqsaaWmDhnotJ+b8PhJFOmNGD3Dc9TUZAPsX6zOEUegr+ubIX
njYoNx2c2F62/RZec3Lz31RQzOGHyTf3Q3tpXB5qeB0JGIN836rT5TZ5Sl/HLt9Ceb8w8vCSg2jM
rE4W9I92JndfaNJP3EJDvk0JIgV5vnI1+OYI+Q8VkhU92FSCxFKwcUauy99vY5IBAyiRzk/HfRsW
msA7n0gXtuMfkY2qTiveeerBgD8ytSw9kjU2W/oxybjYlFB9vRoVDTDu5XG+9JpIvefLStcwOoK6
xPpth/yAG6jxvEM9fhJsl3o0x9hDEN8T0XXP7zE+WT95fQhk3SFsYcTwbeGSXWFX4ZP3wmcTeVSK
h6Rz6UzKf6RXl0/JdI2+ArtEhhZh58imfSvp9ygh7MCnVMTmgAs0ythhb5awf4+qbPhv82aaDp6n
MPvS1bwtEW8ItphggLXokAZ7NE7KCfoLWBO01SgkxvByQh0zyzZ6GRzieeApKVy1EzMu40epIVh/
vIRSjKgNL7AaqZekqP1Lj9usCG5G4oJITEEKXIPbsBm6dlB3Nb8MftsdkEH1KleCzG8p0dZlsWQL
F8+/bccjECT+daYaWy/HhuQ5IPNzmAx2yP5i77Sg7au63NXdRLwcRuNynWvS52UE1md34JpKjcFZ
0VDkdF6VmWh7kcUlqshIpqkjpRtW13SmPdqh/xN3JwPjXJ4MaXw9l/KRTrlSE9K61J5X1Wwq6Fwd
vM+AkRnR7wy6gP2MrvsewDT6sO5T64SWa4MS+jJRuX1tV+xcOLXXPrEMTvIATm1E5/ZQE70Ex1PG
a+IJINvsZpQT1ZjHsVeT16+MR0+cUh1JTXktoQ2EllBynh2IvjythfWXfFHP+8gg37TEBrjFOein
kbF4iQ9o00WN7f0y9srl+pQv4+W3qbhzCny/mMX2uaq8BT5XVyGAE8qQdmNxOwWXejPNl9s7iylO
1w8WHFzvzqDmO0PCGPQOpElz5A6A/tWCG9uGb4G7tJAXJBwd7FbFPMkELsgDTrZXYmBkoX3cKhyj
+hSeIiue7tT3p5IwkZAuJD1bkxmTspN2sRvT//8goOECmHDJp0BxFXkaVbbnPL5Y5stBak8HHEwQ
uiwFMOCjHLoh1HiZv6AhnnrCgyKhhf4Gduwda/URbGfZn28JBChaBI8eiSumJNuiN7JlSkl3qa+K
3J2kbBjXakAKIibFVqyY2rma+1LDLS193ZO+me2dj5OOCDMBhL3KYF8EPWfO1rNCA95zUeelfLec
L1xrOE676OCEh7+FMEu9qDG8dHXvDr6izmDg4o7Y2VSPv9KvXnWsXFIGaXW9wiUyycDmUr38g7Mv
XHATusD0sLkfJDRH8+xOFASkl1iRjSMMu+7iWKEMiAvDc/bnLIDwOZ4vhE+tYgE8AJAV0pD469FO
TlVusRUshu4ZIuTBnRGguwXhwKVOBv/Yqo1XHafbj99mwKWZ2FXPbQhWhYiIH5BxHwPcttWD7wKI
PzMpcJxAg/70vB66xFoMtcsjM67DgfnIWqScbwrP8gXAvr5b/5WHSGyzcfvPd4WpWbX6rhA+d/yt
KxRyAwGXxNCJScuViYMuKO4qHI0QDaCiczj3DMI78+whGLCCa1ol/iHgogFdP2oeWgdwZoOYpa2p
hfmRVmKpRLlVILQLlRXiC1U76u6HOo2z5+q1pBHGX6WAzyVoLHgsGlame5w0DUH44MXmRdMh3sBC
eUtmmLz/J4/PlGJzmIh+lmNLX7t+V7Qc1C1XGQ0lB0wbMLHijLCzNOfGPt0jusZShe9UH9i2VYl1
qchFo/9dEA6+WFpMiHcKgT3c//RrHFCe1qZC6+zIReDnLiKPYWInHJSTPS9GOFYwPM7AQlrUPwMi
iIsWp5CesNF46OhJNh/w69gnwlFWM7SwCoBBzxBdG58tM/1VrVLUw3jIN1zZ6zSuRGyiKB8iF7R9
ZMzYjEsVTZA8WyWnSHgUd8po1tcyTBz+pR+jmHqyx7KD1Pm/zdrMY+aj16EofjKByWsUFL3taaEL
9Lhisd8Bu6LCt/gW7gRg8tw/nw91iEFIXo+217NGdLylh7I8uH+bnzb+nW0IUQOZI50/pOsqdFLI
zt3IxX+ANjsmVCwiJnG1u9SRSKI2fE4yzzfDgDU5ue6WEDpx0L2r6aM5LadRMCXrSJIypMdMSW0t
XsbGL7CM5VwEUfNHTe8vTmAQAtmf6SlJ+njjS/rTz96ZifYVcAG5Vj8xrg0Dt7W+T0R1tduua0x9
tUTm27MWSqF7Vza3ay28cLd2H27xalx3z6ijLXVlSgkTQ0d9nz97LHpNui7ugtqh9eoAMjAw11hl
bE0NLK46zA56E3cYjDkO9LMLfe9bauiKmuO4sR8PBPzYOa63gTHMCuxFfdqmFcjZwYWlfJKfm/LK
iHztDPaRnuug0V8FHZC8mstWCGNs4rLzbx3ZLneCSSU1I/S3cmxsMleQU00wLYYI/bot3xsOE4TK
M36AOZfHW8j3iQbGYpEN/7D/9Qwmg7B7um7S2/Qm6JvZ6MUJTVIvhsHu+Pk7hUsbzGdnPv0RX+wI
ye3yZr+LNFAYxk4CfszsW7bELLoDmn0NCcKjh9vjZOyGvL+yFp5F+LdekT7kTcrrGKckqf6gsyS7
6U3ZDJyEJPBo60GP1DeIxu5AXi4z8hSIwQVcnlrwOh0fNs3C6mnDfkQ4C6/g0eqnAbjgAwBYlVpv
U8erHA1LR3JimplHclWNg5lQkna5ATFw4NBIEvk8QvO98bJKO4tkUqjZbGCDztwLk2CXx9mS6345
kQK4+/+o0/pyr5zxCXLG7G+LaNgFlhjAMkdI/aH4h03hqUvY068589wtZi5CObnP6OCNjTIPXCA6
H4eQfjTiIRYk8F5bH7ImVAaQZhbTKJuSYgKTU8q2PYPu9eLx54nRK+iq+3Qh9qrhDDF9jzfZGPBR
8nw+Nh0F7wV93JXY5LoVHb5nTfAad+0wN4d14nbni8DPmjdQiN7qGNJevbWBapG1E0SRyw6nhS9Z
h6HTKwVikYnVLrklk8TlA6wk9EqzpfrdU+PPaY68/GSn9Kw29pw94So1ubzAY4W0L9jEgeYr0AEp
Sf6uY1sm4R6EFyerReMXeEV2K/2540am3rnSiKymattqwRRfixwWBRkvnsnuKKWbmR2Ki9+f3LeL
G+tAs08Ay/0FaIpTAv4FP7WOXdHscpTfWbJbtGFVuHdXGsh0ZKY2VDfUcsLa3egzpAOp57VMvr1F
LiBZoVwJIPSZKO553hJCJMomNYKZ6o8eTNlSMeBs/QDdvSWuTMkPMG6pmNapVWfLu7g5O0csREqR
IqMlUWOshRHy9KCWWjVaHgpHJBy7ggfBTBf66iyrlIky2faSRfc2IBFmBZuy1RtPnE8u7+/vMHHz
OaS1efBNl2OVOFTmQinbznq7ekyJOSyUPDL1wqszkqKF0n0KIbcBOAr+V+aPHCpkfcG5tz4Y/W1Y
DLjhigHEKN/DoXFgt35DeuuLoy7RvIeRJISJtAGFsWQw0x2ss/oe+KVui1pikOzMD3k8NPmf/R70
nWOdPrzWf9+uMUV2ySzffBisFUbemcXN6zV/K3eGIusk/lustQP7JaS0UXHKgyxjtZiZIamZ/Fn6
T7eGVuAvykrSCDkt/LGsCuQJB9cMXq6BZfRfb39FEFiO001vtbAd5+OEqbhEriMz7xVcMPrlQQMp
HfsJjUeVGnfVETdm0sqR45ylwBNEmAgn8xa9Xyppp9T+2e1XZIEwuW/hmHAJFNkghhM/QHHbz8wt
FMuUtig3X1TJfW24GFSs5YFH9vfl0/CcnUSe88OqVXxmMWO2A6ZnbyzFs7XZ3AzSR7j0bOKbqgGw
Qn0jMF6h0fAl62gkSGT573SoLrV+zbtPj9L3YYY6xoslk/VJfFUiGvAeeVIRSLLfO/cw9wmDJ2AQ
VoimgTmLDHfPDSG6cu6Kzr4Ptadi0OUTJtxEz6JFbaESI35VVeu2awX6WkxrOvNomAiqdBsnYity
Xv34CfUu/HDP+3djnPN3ptMZiatiylEHdZzgGCWB5nAu09a6krlMweXrwWfTW0Mos0sYLuTPg5Gn
jSIfsvx7/UzlGPCSRsOP+8dtzrPMh/nD21nA7EGjXeMcE1jfcP9rYvfJMleGweDIEKfo6EtpocNR
Gjrq2Qsv71ibfW78dKABiZW44N5UkEcd9DC4LUNs8MySSFqizy+3JIVJ2Q5ZRB5zGwOjXb6XvsKc
Q78HYz/Ql7SYXI3rOUM1Ci3SztwCja5bsIfQZC44Vv0DnBxrtXpxfweP4czqJYrt2bSCCrMntHw6
hdXL7Kd25bFlO/YPZN6UttCvpzPGyzCdy/JXGb3JcVb5gAT0n4/WhoEBRkFQ58jy5pqLI13ZgzAr
whT5f6yw7HLs3zkAEzRa3++hgxUhR9RJiHyEyhcZblJexIzYtHWJSIa+yztebnUSdAFIr8OUdpmk
pciwgOOEO/sHFTsnJeBfx5h2KYLvdfD09iXprwRPqNq18OLOxN/93RGLbpUjGJvlf46aqDqZNZXI
urlWbdznA/zXX7UG2/50NgAYFDbl85BYCA0TMHoVyzjPfXI66yUM2Q16DGFbe9l9smwtByjl79Lt
GYUdPj4CjS1oRgHf43qs42eqq0xSrhBHhgUq4K5bg/8xRSiegvosEzzDE0cdXV9w9yPvSvka18gQ
46a2u4TOc5Y+iXbym0sTkmzLh4opN23j+qbZgUB3A408ToZAoroKJMSSYDoIBTk+4bHe0955ywlV
YVxJNod85lJ1o00E7t9kVtaPSZ8ssEOG8fXS6S/NWrIYjI/8+m0ZhWZRWLkqs1pM27MRVZKTsziS
pD/nRIooSooWuUZ6GvesjnY73mJKSbk6qRnchd+pHdHhx0h0QMl/r8NtyFWZOL2zEE0SoP6ZJIxY
SKnlNwR09AzkZE7K0lylIgfxYauO4hvZIY4Zp20XriLIZhuDH1XP0SY7PQo18HzOLwLdfLqmjMBs
SqAumjVLE2425joqG7u29qH2IXyiXMux4HPqzUyxK96JZKMK0rksPiVJzEz2cVVdXfAyDtTfcAfx
Q3OBDEGrx3V+I12JOTMurzBQPKejm45pdAH7J+Scc+ASJvmFNkuDu9VTHZyn7J86KWD4Ae7f/OsC
1SzWA5jOboBUveT16Nm2SR/q0PhSuagLfekHZvoBknWrvvQcthNPlH5m4hEXC/CKlCcrjfzrF82E
6niyCFTC5sh9Bllba4WIXOg6PELJA/+BTVDYZrQuNFYhUzVtlbhHmhyp29OiM0m9vdQs1bKgpvIX
RFm/1vbbTxAmF9MU5O7V3/Ok9ebU+MM1ulS5zGXAPtq4IzpUAboanCXL3UuQcwemPCchp5oSoCDN
DNS0kI+0LbEZwM6MWXJ9Te0UUQxti7s1aSjAoWCKyo8vsOVprvq9KptbWoVIN7ebRQV1lzsi+Nqh
I0wgSBK9ntMr4eypEF1NbkLjc6/3KcVFhpjYq77hkaXlK3RHJ5QhuiihwWqaUkK0jg62Kb1ZwbFt
v2OODKpZak968ooZ3SIfh6rnLXlG2tIedVk0Qo8ZQjlPhLDNYOudtb3j4tAzCF1GtjHgPhZxbfV9
FgAnshd3ffoHSV4CSnVUiXZdmCSuqTrU71q3M+y0BobCeKv9RgDGyIvbksPFgEkLrEox/gLIOg4f
J+8Xrboye6tsWdl4x/Jh7oWqfoNScR5VWCYD2vURo8sXiJcoyeNLc4l+n7186SxrIKtlUOes9GR0
0fMJI3kGig/hgTqKkD3zD/I4HUGCijVEUJDiU8a9S9JBN3uEmbbkVeueL6s+H5CRo8YG6oOsT2rO
mhIPXl9hKOV0q//GCmEoadhnsFmpc8yN0cR0PnabWoicqEASqs5nb1Ct8S+xDsOMvRGmxzFK6ynh
kdxxpSGy9OnIPKUxGztpwO6/FUN8MCpdd6+Ewm7Ocy/Ibk2un6qHtPbouHPHRF36froyqTiAlIOS
xGyqPZJjFv2u0daRhPDqKLXdDVmkBVupjQbtSqj7HTGIthZ8X2Q+j3rAJxMNcSP0u5yURqpYO4By
/H2njIoyvf96VJ8A6h/M8bGK8WBC89xpY5YnJWsRluZoelECiQ/KmgONpxz6J2O6A5G3LKJkc38y
wt4HdmgX/F+Wul8Kw4a4RJLQZaLvSqQ2nFAtayw2kXzqvuI7KyVltkuCspk/5bdNBCezCkE3nDc/
EdvDT6gdj5n3YjJVE49hX/vivDOfT37LfzJK7MwL4RZn2i4kJXyeYpqiEWu9IX2vhNd4dhYaBjYa
KO3DEhrSdhVDlNRLEnDoMuwH5qIQruzjyWgn6Tr6NZDOQNkYPn9Rre7zmuoOA27Dy6/R59OmDkwG
cfyMI3C5ZxilKFex+yJZkUFxYft9ylwAJyblmalMkmFXHlH0abjm7Cm4FyEtSRDSKcKRZxLsnkpk
6ePAtwzWnLUZDmoD2z+wtzQVFp2iwSlB5kxyw4rtuH/vwtf9c4Re7pbXE9Ja3BtfFaEcByPhrycY
r+WKr9EI9oxiKAigtwFpw3EiUE35pPbNJyMe0w637jriC4uTed1ezrBGWhS/7mtKo9yjjHteQUyJ
AuhS19FE7jI3iDhQ9ZSfSt7FzDyvWR1YXjJaqucyMCJakFRVwzTiIfBK9TITKW+9TocEQVcvYrij
BCZ0y7GHFJjUDXexTfXP8Cmxfxa9Em/BwZ1LcHfG2+UM6jPV1dbkRe8kk6BNv3+1uo3WXO0w6dek
2+i+6HO3azjuzg9JTEAI1HLHYL7ZPsqrgu3Nxy4uRUIwTMOV4LsSRlBF4OQlHFZxBz9zAq93ZjdG
ztY4QOAFTOhIZ7tjyZORTOpx2xV6YnVil6WkUrkIwKp0SAP00bM90Udg1a9CR5HWyK1QGiEvLA1M
Tq0reMJWb1LnAnU8CkHBaZEfURtSLJS3yiHAmkLgNYGDwcaW3c9qbCcdhCjdwwLtGFL323/wW5Jk
qjjY6YzzjqAWlwYhfJosYbwoCn4wGbKjWdVIB7LLr+dNUc3vaeECJThXjGHdcs+w2vlQMpf791Ju
poLiUDWfABnRIosanGfLNBrg1CMHQkZQwyfNLj4/79iyWWfxOlgXMu6VjOY33Ag/z3KUEDT+FuOP
FkK5+EiMjkTvV/VbfXtfELz4p8xicwWMqZdPI8zyVztJ0Jxfch7RFngZq7YvF2w3fcSq0l4wI7Uw
iQhVhBSCkf/JUeh51FQYaGUqnMrLCK9l+zbkUpF2EpZ8wnbh9RdqPLHFuz8fAXUhlmZdXDHbDGej
EHuI4pqNF5+5cGY7ZAvvQp09ZWI/VdcagRnRkqMsoonMbBBVOLa6qgWhyfNM1L+F449LqOhmjPt8
uqUy87nXdHh4jZW6YSBSTZR0GVLML2rcOZyS6QdFPx8hxX9WDUh1GK55E8iv2jKSquT7UqX3HoFc
Qebo6wLxVd9qAsIbxhg/xWq3QOkECUwJuEvRDZ4jBN5u+hnhpRDKrGE8Id3eNzdzXoROZOLq91TK
X6WDMVErW5ro2Yh2/eu9LTEx9eBgylApvIqpLwmi8OW+RLqgMtK0KrVYewI1TXW6fO0sXHkd25kK
YgE2dOIWzk195ihMNdV74WpZEALtsu/8bNHm3PgJaYr2EOiDi9rDUoryXP5NWDr06i/7pjXzHLpr
lBBwR8WQVRXFk6D/UeCFrwKEmHCxeJVTDJsxlpZLuDgxl1tH97Fn3Oz72JFXgdKv6RSWxsGDiCD+
wlqK+aqUMsMYLuVPpNBlExU8vXCKK8Y1FC4bDYrTbilJqEPI+qx3NsW9hK297Z0bV6XABUuGhubZ
qfKvq1mBrP5ircM4cuX1a94ryEkADLzpuNW5yuFBcy6KPyO/gXioDquniyJN/3CDdplND4b6EtXD
vLvJ2+uhZCxBU4BDBR8LvfGQT/06+bMElPYXW8GKkmMZJdDrSJxxCEiY3MUtZWAOANIfQpUBPhvn
qgbCYpAUp3A0NseBvWaIArKqDVI+KgP7pcXRadC+qF+NYm/xp8Xy0KQVCd7M0S1b93oZlYGKCABL
46Oh/EzjvXYRWuX4QwQ9VVDQaoUSBjsWDvF8JnbUf4Qh6UuBPbJBgV0Hlh7Ffa0fY/wkqtE6sbY1
97zTxfIPv3hICFeYKN3tt24jFyJc4SFWFdXeCvp7Snif5lfdJODJw3a9BUMYqXmXCbudaS++F9Ca
4tdj4NcTlMoneqBuS16ciEoZItdXHFdKnfQ5x6fiWpkWKFE2k9UJRd6dvOhP8TCmf2DtmtnNwycA
XLrbKzw/urbDyoGMELx/Nj1jQMbNz2PUlfz77vkbFH9YZNFj1qpOLisqzin93n9U8Kk5CCZKKR4b
jgQr6TlUlc9E/0djUfkR7b68SBYIYssycQEEltElzl7AbNX9ko73+ODMgncSL//MgJdIZduFL4Tg
TSWf9MFZYlM55VjlkMBVPCXwIOMbhnZtjspMQ4rrDRB8DqZEEcwwXvVjgtFLXrIhMfg0CfJLjaAv
CW89/nl/NbUVAloUkZxNLrzybOBx95ujIBNhsl4dnnbnQNSS/N3EuE/Q8XiSzizfwdM5nX6PXj2D
EZzw3Vqobi6bpmpVH68Ocx+Xq5UY93WHEBYgHqEdpUjvPpJKyS1hKLopvTeVa9O2EtxdjLx85szi
Vu89M0m75Spffqh88V+cSX+jOhJLtxh6TQHkG2qQbmPESCIHC5pCwSP9nWhkkb0voKqRP2fMYm6F
URE8OW3zU+CCVT2yTnXXm44nKZSAOMB5MTQcduNYrBvEPaZ2olQNipyyeF8cBk6rlg8g1/HHV6kd
bvYQDCbIs6gL92XzD8319FEmJAFFUYOimozro3m2x4XcL0KgQJngrcqcjV/lnp36TI1Os7Np8xDH
61FYSJupOFOBkxhCegvHbqRwjOsot6QvArHOajQYQ+ZXeLZXR9MCI7i+mdjHIwFi+p7iM/nkN8ux
H+jEzfWpxJWrkALNbPYV0IJ/58qocLefuDrFqTBrrpygTbbiyJCvPOPhZgf6LpJdQeZ6iI3hWSSx
gEB792/GnuwEpLbXgzDux/21bl4xX1kGmqhcuP/7hgF7FFcDqHJv3XJTTjvvuuVTqD/vrNlDSGwF
+4utmSWeX1LENums35Eve7TDL9xobvOVtdoljPp9Hq4isagzDpU1piRmeYl3tUsV1zExzCq1q6EQ
KkiftdJI0uGVKxnuQh12wLs4pL2V3r3tt5+lvHcaaEnN7pPJrWC+Ep12LG4Gxj7627KluF+Sz990
SRWnnJvC51jd0tWSWnfPS6zlXHrjUdVzEka8naYMZWWJONfLYegP30Y043MIZW621N4U5b7C0KfR
7BXR3trJKeKv4iEfm+eIQInSdiLpO9Bti/7GY+m37ZkLsFf9fLKayTVL3lPgXervERPBgpUmR/re
1NkZZ9xBMTsf0I0LDNEz8zCTQXytsaFHXb/bkYPqthCWcObTgCAvcIkMzLUhNHFPezx94GbWgYg0
CopZcKgSGm2dWveu1mPcKc8XD37G8FCArQpsbcnVON8uJpP871jTQ76GzGVxrP/qq7PsQQjpSbOZ
yUzMpmoNjFzfeZ7vC5uz4GHs0rL+tJGIkR7k6M9oW0QvHXiIM2atr/uk/IoYTs+2rBWQQjoknc6m
YaFwRPRl1aaQXghi3FScsMDJo0A0OTQ6/hsG4OQSwVH/CnxFWxmd7hNs8ClCtWivfJPOrvDA8699
Aca7eA/St/uh8AZkTZFBVawh0nxWtlyaG4oBtEGpxIjiFAehniKUBKZzY+WIuivaVF9yAd7cgiIY
uRx0VA925aPJcDJW4frfPTaOICnf6wBQ44aGT2u/PqlcH+T1MAhLKMRF93Rkn6k9DxQaeKj2da1Z
e+dEuA3MjqGSGVCg6MRDwIeHhCiAPyHyeGbEfovWuHbP6KrAwv1Wc4B3KIxSEGbrM5D0MNud7nq9
K/uvbGQUktIqNTAXs0T+TYkvgBiZu9zO9pgekKx2SYrENoRzqc8bd4PX9Q86ngvoGtaWT+zpT7jl
6NkjgnsJD803ahLFG2oqjmeIz8Meo6iQGUCZJZXFfqunF/Spq8qd3TLB+7JHOKvcC+Q0DEP1105u
bwYgPOG0ww4RVHSwvXetKwayiGwaLtJZ6neVp+q86eIXPfw4oq8iJ0R9HPIwfZuD/qrDWJZ8JYIu
LWzUUFrS2M/9QlUyZxdRYGTkFkpdvbjKR2JleAt4YDTdyr836obluv1QmyJHy3C1Gx58T2JO5ErS
CrF7ZxA4bOYeq3XggTxN/JNlS3GmPCKv8rA7o3ycrVpOPuEX8BQVgwooHlLkMfbsfbf8GOp8mb3a
1e1J6DAvZSZl9+X/CinUTunkqxa+YmkfHf672zfAL4L53cNA9YxXwQ2dumDqvF2TYznY8x1UpjiF
NiGpKCpMNh8HqXyUObdIAvmo0Uluy+jPaEFYedmrQGCz34xJeTU0QO6mGdC1/dEGVv79R2rJUSrO
ZPno/mHHkUCm1xASVocIE+fdcGXUJIhIPykjgv2+MmkNjnPtv/oZvKzeT802lLuHxe6AgOXqwxxo
VdJT/2sMdAPKtl3bknf4zZEqax1SyHDtNpLEj/eGvoXoyvLtFxpHfseyo3C28OnXxMB+/GeXtWXm
UvCGJPLXoa0t5PYkg1LNqMvxzlWt0zBSaeLz2pfEvPSkKXFel3to5anPAPDQhBkTOPDj1doMqcYq
30nb1zmJGyfkI4TsLoIG896U73MISixeRZJ+XQcL6SlNjuapPGxl1zY+MnQGwnAaDifCpNM5wv7m
pYfYFW91RWbqYK8OrdDnr7nojCAt/N8r5wqNm7cibybg8mgGz1iADV9VUXkiRK8hvlk7NruQIkJE
FOyNib0BnCltIrRKtOAoruHasY4LKD+QIxZefpK+9LB1fRadqQZzdf/Eh59qkL4639bEiwUvdBeS
yc/ZQMlWRTGUo8q/r2v/XLE91Cv5oXkNkxB7PY7pDPdjAfigQxWKmecEfwdOr2ANPUDiYE/L1MXv
LgwuqwJZQDjtPVVsMam8zHDmBALCi7X+TkJuvU2ABw1MnQhZdvCkR78P5Ep3OSgtK13OBvsLYmxE
591gl80Gyhb2XBxgmzgSZ+IlVodF4jSDF3wFy1uo2+iTltyUnFFcrxYYf0V8U6t510aBVKfRJAeH
NGGXBmp6bMgc7QyDBpS61C2jRzcbiMq0Phi8nOg4IrvHlFdhsZv+DkasIEUZ81lpTj6NN3DwDght
yLngUSx+zF28CDvZb8dWhMoaEIxxhQE4Q+/0tEjuZOE3JVU62PHyR0yGzqQLzyk/fi3iFsZgRgu/
nobPTuLNI/Vz2mCYFRPKl728qTMdYqv730jugNavYbOr1timVz1nUfFvVyoue1wCwYIs2N1gZ3gk
IvRD4JsqcREm7LR1cg+rAq5hv6wuGz0Iz2TMSV6gv/CbzP98gS98IpVwvfvMFpKJz4flFY5CaZxH
sI62tnIhGvMXEgrCCR+a2+VodDE/7E5eD8ipecFM0MkCv7gUXd9h0hS0hBvfQYoCnWig4ZDPWMXd
aDQqIgXxBV/ffEjOMjM9RbQXVeCPVLT5Jt7j0U/77D6sNwRR+hoqRFsrTNUP4h09qqtsfDi2USRV
MKWOagVhQDRD9L+7l+2flM+bX1bQHjJPLuRMxoYwDGBjeHnkFQXqRWdSgnv5PBZiQNTCiS4w2PlX
/U1W1vzB31xFtEWkFWAPNPiofklwoSTLWIlaNqaG40CJW2SoNPdqUXgTnPwCoZLZjoZdM/0Lx1qE
xjv4H23pjMr/VJHKOuVIjhIRva4jJaSvi0w7SULtafhrfgbG7TyTY+k0o8doG5j7hBDroZChz69m
Wj8zCgmMnafzx6cp9UXFm0Cq7ro/w/UMH6ysTLSBZENPjk6lvy3yhrFBmFfw/ComdXmU4QIw1xtA
/0mHR3D2cWnuVn7j1DcieuwyagSj6qpe3b5u2QJlOnhZ94PcRhDNiibvBmqGRrCt5EzquTBQGRNB
fcajSOdXBuKvABMfizptClcurK535TZTUpV3ltu8POmGCJOkIGY48INRijg1lXK+L584RZhUkgd2
9H/29Oe9BU4cktWClFSmDjMJ0jWM9kSjjV+pg0TK/vO6jvKtYE4VtnQR5RZZjPEAKR4jk6B6XPHC
0Gla1Ccm0UOUxXR73dDbqivM1hp/UuOyaBg6u4AsYeMr7hGvFksEJt8V7HnNy92zUnBa6MYLgByo
5BKdzVOY4Zfdac43l+b/C9ctU5TX5gPWlGHGnuUNVfO05pkle7MoEGBFA5S9aR0qsF4h7SIlR/zW
WN30eVYU1bKV+6M8gV7u+CCGoNcnaWp6MdGhqNXmOnesX6zW0XaWhWsL11xb18nGfhb6S74vz9Jj
2IGAt1lEFFShY8l6h03wFh+uo73lTOsgK+oSHPOSPErQX7RZq6YqM/tLC2RSxRfm8hFDnhv7Tu02
tOMLY6s3BJA/2lX58oOBajbtkQ3SDWN2m8YBIK2d0jRX790iHiuz7Iqdb2b6iip/3f4hrxg18U5w
K5Ihm9oiVLuuifMgUQKZvlOccI34P5SaQWd3/y5Si19p57ToHwKbJ+OMmJidXyZbPBxzC2EEmpmG
UMh88ozEvZG8Ivr+9mjgLqGLZm+haLG5mdLoDSHGbL9Fx9Q1M4Jf50s6HDNMSNS+Gxp/NP1actie
c/1ou1P8NwZmcpPip2blJTvKBntcr0NOr1dGt6Ucl1zHbek9f6EI3bwrh7tu1JZHacDBoYOPBDrB
ZyhFFV045KXerlHLgt6h4NH12GfY2ubcn1h+wjb375X5QL99zfFXYt3060zBDWiNvbNeKXVOe+sy
RcJABZab8ExQFywCFpi5sYWtSrVb5palmp/rO5q7ni68Xy8li0xyIGiNuqSqGcgGtLxTY8o3P399
gNLPRm6mN1sf36IZbwRTcmhXTvBNJRzfDhcZLzVJUCToY0LJELc7xqOA75FHOTQrHSffbQsoHrnf
3+i7VhUMF4HUfaoYLEJ1KcYi9gXBRRmRx1/wVZfl16PCqt8hICxCDQMXo6QPtxHDsyQFcgkmparY
tO8KzMon3F6iBeihNCkyrrfyjTB57XDEAq5L6u/S6o776ASH/DV9jO4es3/M4328SSC7zBDgt6Lg
fkHSKiAYchHUg3R0MwApVXMnWhkpNevgJSSa8SSyhM2ZtFBw39ZUyQn6+eGCWxLKjDAYrglzr3Xc
hneGcQjXtc67KXbcQQtS8HDDbdB2LYbOCjyDjpPY2oEHAxIw+NQqGTnreIImX6+D/0WDtR1y6wbN
Wrd5Y++mehMj2GXYNBrtA1HfFwUK+fwgAuQlG7G2p7jECYVPCddfgq8bMT6wWYEFQljFbKnVkc2X
ITSaeCYPanNlZBWHaey7A+9CLonW2Ij25pgNJFsMRO1Z4+ahkxPqiLPeU5gGK9dz9+pcpJW2yI6n
Oxz5D7E4k+5NItM/Q5COWF1FsyvSM2Q2Q7ShkcXVzjqoPjNe3NBLXDUhEos0hzz5VJeaMJHqWx8l
OsAMpBJu3L+gYLiYbFQKzqtTuRlCnQVFvi+ZCF388s6OO3r3tT4ZRnR82ZttEVTDYgbZHerTjt1h
2UHyWFrurQWqzn/Gplod199EHtkrasSa6dcF6irMlMmCx1DY4kUFuv45A9qryYliRWb5eVbGMjs2
wU9b6iUeq62SqnXN/VwIq8XFX8hgxZkXmvknXAwtv3fIUk3sXLRdJOX6dakahB/HVw/xi3rJy+iN
u5U0fSMQBgqg7hKyz5sToPjfIOkAyrak0IEgba2vVcpRLQZtNwqWGOEUn6EkNBwF9+25rpotMFRg
WI51XwsJvvLzt0r8jCvVFeeHRTcOHjvv0Y/0sHNsBXa9arzhUVkkfN6i7SxU1VYklFP9wIW1V0dL
rcs3l8hRKZsYuiyVZqC7LSxrM+OeQXXWZRU+Z5j+6/8eSjzKh+/uhyPK7b7F+fZxn2EUylDm9i7r
hEtGHvy2jsfmEFZ84IW21CIJniw57J8GFCMstXsJyTSVaQDkQQoO90El/GzYozUhA1xDDcQTF8dJ
2+sEY7SbVquDoQBxJDkX3ADgTwgfjtazdNbtVm0ia7vt7pZxTo4bA5ewzwpLCE9mS2uCahCbBWiG
8mixZeI1Yagdp+0q5OeQ9wIrcW9XtAGGVtTmmaCCQLc9wkQEmeSYvg6nTrnGaVyByJVIRJeNIeWK
A2+PYVhBuLQScmZiowVRqSdoj5gU4UBqMtQV9EhEfxAKiEQ8w+Xa2hkqv057vr6yP1LOl/LFKlH4
id3PBs9WasiKSAbOevabZzf1d8c+oCkRofCMl9foVc/BWXEq9yAnSC6TH+cHXoxdS2jp6SwWIppi
dUOZIupm955e5WWFLwlemABTRt1fxB7J8KcXYT/iAN5WUaDBw/kUz9USZKhR4lRHLKN9cUQbrLM4
cxmXn4ysZqlFXSYQfzwWQL95cIn4sBJlpQCSvqf7O5XEz2K3mY6nv3t8fYcnbwGudzsmNST1S3X9
pIk5WgabtDGnSN8NmA2pyYWBuT9BU42reV0m1vwZCfEcdZaw5HGuksvvUnxK+7jlom82aAjK26GG
zIuU7fQ21UUWGIyjT+l2KT/QAdWFmaMFP/93P3UbxMXtiUcIz/eSsns6FtjMkkXxHtnEw/COz63c
qbXo+INSunWuAP+VxQfHEDybRWVoLPLAcn9xDJYeCEUbltKiqsN8XPTEHAH/ujjPUnm8Nw3AK+8A
ll8J1leyaR9tPVnua9M5gWUAKGVd2Lpl6SYqMoiG79fspoEhFBBXJyZJ/hAEK3H3V4HgwzZfUHv/
8qnnhp974WstTB66fBNF2Y4wGh8fjnRcAHR+Wi8Z5kEgwOu+tZQyLUNXJyAi9y7VqyEx4L87cZaS
GZhU7QW031SYMItnYbVkS5gH3VeTlI4AJ7BGphk+0V6Ib6XLxJnD4T8Fl8BBnMZ9ZsCUFw5R3MAG
2gqz8l7b6skDsR7UYuvnqYJVihblNXPGN60yUiEMs3Ks3RAIHgld4TIYh+4LefzlwVCqlowRKB4L
LYNE3vbYKj8zxte47wAHr2mu/Jm1yVK735QotPgY6hdfXpnxmCDkHpKZdjkmMCsnqzbePXwiUxhB
Pi2zLWPBmYfEi3CKcQRs09qxudmPKOg4qMLsrTh+5g9l5TNztoFqWpn4fiW9ED28cE2CWqj5uAGZ
pI8tXrahbZsgiK0pOjnvShHK2UZ9aaIMRL+omBNb7bx0fORWIMCielR6sEBSpt07pVGMWxxMMHqd
bX6rmaTO/6r/LET0MjgBYfvBIZw6Uxyh3PkrIqkeSsodF/6a2QDyAm9NXpXSWjv+d7ULK9I9BBd1
wI040m7ZMp5vPhQpkwz5LqyW+sD83oqz9kB4843ljNQiz6dXaTyvOFCSE0MZuYrJdh26dbFZq/fm
qcOBxEfVJ+e2cbG17xGmW3fmMcmw5MLW7f/E2ZmNN5CbVT5YzhS2BrOHBW4y/U4RZQdMES4X4uak
q5mRfMW0ZqtKGYL/hXpyKYP70pa2t04SB5cl4eIJY1YWkMz09fdcPzdtaVeBrDhz2a8xl+jZAgrY
21OwMp5hnfwhVnJbwAJRSAN4oyIcS5Vl3scl5jt1rAja6dSq2u/CfUYQAJU1cufTfXn6AsU+iI9U
7e5kmSPc1GngkZavUtfVfmvLUfXCvsG0rF5ZEV3BMBHHQbytCNgBn+bgpVdB2RXhd9l204LEH27u
sc33Jf58UfaiXIzxMpPUHplBIv+Eo2E2ipL6Gl1JM4PetuJAcyKbC47VmVNDETJFZzbDP/L1buwT
v41izX/iVjjfhKOWBGlEgH8WSOwvMkXX9kP73dkZe9vT2DnDhAcnuOg9Dgp49IveOrMk6QDuytjL
JEH3DA7wV0oGiLQER6jmuK5jVQPz/GyLLwobRSKsPFJRV09Ht5DZRrp5MN9urIaXGKtJ5/VYeMrc
yHiUAbObOifXclmQl2+v7xK7pFjSjhGs/nLXJAyjAgSe5bxfd7hSU7SbLF7on2Rj+faJemIrUWVC
zFNLrYh/w2lWeJP9fmq623TBlpl3RXUjvkz5NnzakK5bipOZ45wPaX8aWR7tDU9ODcLwqdCtb2ZO
IEdPlUi0NxePvgN59E7BasodlAwge81GtgYvwtwBu8tMFeLqt47z89qU+ZUUBIyBsy9cz/CfjjRY
AT9bWIrKrJ5HNr2GQ/uv1/E7hpu3ioraDOL25+lND7u0zg6NOraOuFxT8F0MYplVw5/Z8ZNlr2pT
gTBjfgngYSGxeLlfSjCWBG+9zYmvVMZNxaAoJDiUL4ySkhEjo/k+WCSaUAAOqxncq62fps29ji8T
ibqhAFr8wjOwPv+3yj6W7DVa8O9P3Y6w9gWYz6FD4t0paSucxu0+hOLB17AExD2pA9+VEkA7H6ji
IKzdar8WVYt8j20RC4xSRNQ3xRE2XOrSywJDGqvsMsSYLdPXwIAAQMkdcI67T+Gb9z7NYV7iW3AQ
tpqcVHfxRVY7GnNjQonVJNwt0aBLunaP4QEOuDwsJ3zRwotSKCCitFI1PS354H+pYdKiTzlYsMIW
oJddGXy3k1opPthvbwf6c/DqkKVwF+x2BRyBgqFDcmUxCXwSt735q9L3IgfZ2NyLfif4aS2+/3w3
hKiL+F/5x1GlH7Ov4oOsfVz9KJ30VK1/iU7avfcuLN5SXC0kEA5ubGo2NWuejbGwZWygxbtGP/oy
0I2m3bEtuJiAUNjHjspLHI4cEVOkDkhEzZGXXNsxd8u1LiwvIs94MalmDbKFcdHZYzbx1/p/RSo0
4O8QGfagN7YSNhtAfhtvkD44BConRnllRKnd2CaHzFxH8aUVscsZ81G2Z0cuJNT8pCzgVPKl/bkl
0cWEUPGkCnj9qeOKmsnbqu7VY5xcPo7iqQMTwW/H/SnG/avI1n84PJfx+2KYmTQkmw2a0Yp4YIb5
xdjGPmS6E2QKYspWFqjO/vcAKa83eprF1oDMqlPldOntwgUfGSf4wAQAy+dVgEbY4mL21DAwTKid
u8Zfx+nA/oDxc/JIL36gAN/oc3v/P6wy75fjvrMVbaq3LvCsCU/CaH4SjsI0MR306FHgR47/DV4h
z9W8pUsGwI6b0IV3dSOhvRI+vuzoMf9owu/+nzT2R6QKHJ4t2IVpk04d8igPEbc4OPpXVVSLGVXN
WABs8mdMCSp5tgyY5EMpSCFen4Q58nLhKYM+QKTyVjxp97OZgngNX1IwdvLckNWIFtbWMMlaXT2G
L/FGQgzmn7u32GYcOxCKxGjZGiUgdHhl93z54LP/iz+KsYTeK6Ltiredi7caiJqwRbV45nUNrESt
Fn3yB/uDFMKLUQNIE5IopC5Bk1xYzesIprqx88VIg8FYx0M9rpnN6UMrF5G1KocYushXXbGrtVD3
MtWqg2J8xrvgY+dQ91i+FbhAuJ+fZnoKNalpz9FaPZwDT5s33WV6gNRZTcF49OI+01pRdepIHW8P
FY2+6gr8yvirPt1I26ctIeDz72KDS3rpppRUbQEu6nvuu1a+eC8eM4bS4MGl1+45y5Jr/n3kDI6Q
5rFT6hQubWXL+Ju248GEF/JyXM1TZwhBmyMhDwpeJPIbekl8PNgNB+ZiVygnczxwN/fRLenNwg9y
f0z8lbCOXXpzHoGZrLBIjaA2LCVKOFXxaRDWU5T7Wn/s9UOBx4EljfB5oTV0+WwWOsIp8HT+UWan
lem2Q/ae4ejdmAYFVP1KeRp/1l27l1jwTp3j4mAhVsKiJoqYDOWKrua7hJKZ2NwMN+A39KrBb41I
KBa6evwx5G8SOeqtPaCDL9Blnff0ccVoda2kItkJp4RMq+xPrZgoc/wWz0DuKypFYJkzcLf+M7tt
94IAqikSCm+ezjSFX2eNDj1kbutmQyAJ9yFYL2P4+Dj8JQzherHHHMsvTB84fDaybZEZ9ultMMPg
nBOc8TVygupokEy2bZFidEGZu7C++uRDrws0QNeP2UBiaS6Snvy3nIyyGAjqknw5/g3OwfsVq5SS
8uAYQsoMVD1w7R3NFt4JEPaEONHz6gT1K/k63+i6HrscOCqAFFL+UFCvIRaW1e++dO01HNur9OJA
McQwzZamFdeiIgv4kGyN5Qi3dpg2ly9aHHjaZl/eJk6jSZ6FjGxGC6/k6nQfjyUTDp1h2UeI3yOy
G4DZxvxpIxiGkdFI48+uPmyf5bRFOsWgEW/q14IjjdOejSMDEPUAVkFZe8MZrybhkMgPt0/QvigI
q2p9pzzMYdEOjHsYcFVbqH+K5Jf09ty9P5sEH4CKhyBgarfgCk4XDXPNzpDT/SKg2tjXjW69lzmE
CCQ7CC2HDdQU09OVaFqPw11Kk74wge6k602kZUoxkund5UfoIwoDLs36AKtx/Va0iwIsmJ6ikoKD
HBCSTqblM/b8enLvQWircjwF5NgT0RuPMhKVQazDncYmyvJh9I0qG5gaXF5LasSFFdkZd1YSNoO4
38GKxHywMLeyFOAlszIm3/6iDUxWaP723IRH59cZXSNrH96cA3QMOSOh1thqEbJJAMHWt3EjWjMS
aWpHAh9zdejDr8KlphoOe5IY/WvtIF21QccmyPqgIzPDW6/X/HZsgW+KhzIXE+HQHEH9Z7cwS7er
o3D3jP7Trm1keN7lgIzSXwMud0Qrd4adUoPd0uGJkUyqZqHjeYjSUskN86kjPW0IqtcMx03Vqvam
Kg6rwlsshZ0JIbZc378PXwk3voNODiQhLzK+JpC+3gazQaOUIuvRNHX7gCElxgdw7rzMvjBe0LyS
+zgra2d1vdTmkJFfo4wcIqGS/iqLJql7PM9H3OUPIQQjp0gPXl4AIAyIuaEFmZyCmRfR2ZtV0Ibd
aqHB1ILC74tS6Wnv3VreMmry0u7Imcd2cXSFRPVvGYojUBRUjaZNeqnCR/ekA6DHHfdvrCblQ3Mx
Zu1GZSqCciD/kVEH7tLslxXXLd4qAKxIpcNeXrIkjx9jB4cxBFI7AGFLaQRCvHjmxzednKMcZkpB
p9+iJBoizawAySC8ItMJ4fbraXvSgbmLrXfWyd0V5x1mOUQuax6hOKxiq1XcwoKxjpQ9NzN1BFVH
NmeqyqJplELcbQjFcaquyXYRxfACeg+uDZvBgoro9nUp34IGdFA16LT0qS/JzhrHpCofiOfKu2Xg
IPnrhsoQonLbJUdLZFn5Nj3kcXQ/rU4uqqohhgW6Kx4glJWV0Hrmf2A7z9emmNRffme1SerEVbwr
5LV+13tk5SoNCDiofJfxlDuYIMdo+ZbFay3Tlzz395x3ntQ4n4IzlYmfmlS5WJgo/ucoyX+bFpXo
iPFh/26rVrMpUiQawnMy4Sd5lNLYYxQF8wtV93xzhuouPJjkm9Hwzrlct9053a7MFLuJmQmtj/Ny
Hm4aHzZvjbZKG6D/7J9R2T0YBuOqEZAEyrc2f3Qx6FpT4yeQDMp8TBcviiz3fpBAavX8XJDH+2bU
7gCHlEjE0Eg7VL9PsUZ3pfrpIwNU1sZ0LAsqHiPgXo2aeow83FsDJE2i7LhDE6/wn5UvX8rQrdiJ
jYIbe008xJcAdYSgnHKW9nsLOr0eYp+dBYgtJ2G3Q5HdmvcHPOG8GnC5XM6DG5u2aTvhxaONbiaU
H19QDohxQuQ2B6h1Hsy7V92YHrAnTuoqdMaN5QdAcqAqegSeam3X/OF2qjm5I5J2UHzCJ20YXQ6K
P2JFMW/uF8DwfV5L7E10Skh7uyhiUkBTvZ4CkypvDx/wu7m522WGdI7d+vVM2FsTIEOUL+9YFfd1
CzNRRjYdeIzOrOizoUIClTEELUO4IhnfNLyFCAn53zPCL66EjRCf1Kam3yYKqW1if8gl/w0yr8xt
zIz1dZUi1JOIIr5RhiCyOxXrYSOO/JTy9oTITQ7ntEo5ZRK51V2nFQgmEvkwz/C5Uh49/BZVgwLB
KOHEdVoTcsmAiHhAFa33i2kVjkuXZZp1Zh/6fLB/uhAG2cv8f4/PrT1KQQ9nFmVL/v/M+pwa2kmx
3GWSIm8sPbxadmaLlQiueB6jEhdSGyoqTxlCt+s3EXs9H7uYVg9joMURsc47aGiy009xa7zYVVEX
EDF7FRQpF4oyOu0H5i7EfUKIL3+5wZMuHRkVUMMy7T/JWMomPHLT4kpuCcMXEsKt1+zsiBLPBa5W
DE/psIr/sVL1mj+bmifsBU/BiiE3aAl03S3ASP6hET9z7E8Nl8IfMIfDADMNYwCem7iQG24JVVx0
plb0FQ7qJw5RV2FVp1NiBe9HgbQwmjU/YP0hczm7GTrCd9l/76XkJ2JKMkMxypHPKcvUtvbCT+5E
J5kwxCQF1hLp7mJrkNLw9RlUvfQ0ZLdOtSS5DDoN/2PhUD/ohWariNvIKTQ6W0kcCiCgpwWeZ5pi
BM9HGsHc3aaenFzUww6HQw0flpOM1I2ehbyjJxFIA/X+qrGprfR44YhmKF74YDVK8EHWUFmN5lu4
kmRvjLFQrC3IKl4BNZbjzjdAzkOmAne9QSfmhuk7hALqYsx54Qa2WSsDOsomYBMjjBZ94HDKJTW3
o4R5JfyuuMDF/3vwBQBE++NpWRI3BYm+gwRe0pjqhWVGxxDB+CK56ZWyYzDWzseIn8Bcb4VII//Z
Uz5xanW4YbjaMiElsFoWDcm6uDlgYjKw26KzV0/pTTp+2lC2Ty4jcsp9HyS1bzFSQagi0T4O5cTQ
OWE8zjRXn11xvGkLbeeQke7kQOyt7S5qCjCxwNIdIEOAtJCjQ4w+L8pIVQ7Q5MSYt/7s20f6vgNZ
crE2gNGpxdUm52HR4tvDSOLZ1Mc4oIZ6oYncVx80e20s6n49W9hdxzLQA0AGSZSVmKi9FZXPjwr8
lYsPI+/mOPnQCQT+oKF0HrrjqktyMggJSMihdsO/sNXYHKqm+FlLwzOs85AkB0QWvex9kQMJgbuC
e7DfQ2IzkIdctVE4xNqm/P/1in/29oFYx89R/cedD4HQ7Q5zJakIG7yoV2qAsLqks68vrAnRJ/EV
k4ZW1CMRml+QuhjemU5FubtWQdlE5AqGjt82SpOUrd3WqiuvXvJgWraZsab0rl60p/o7a98sIJAe
sl9VgotKPnIXy2hLxIvPR6icJicZQH/NAf2grK2TXHokWAzj6eVFkAquqT6yhFvQUZe9/2iBN7n5
iLlPGdkqNjEz0z42KFIDaxr75O28lxuxsP8RDAS13gRVVSbsvIQ9VKfgw1fLVlzla2pjKmF92IcI
Mx3KcBehwwr1/LANOulb/lO6Gu2gxXJYO9x3T3pClRNRQ0fIBubIfRMQM+grUKdLwntmlFWldUcf
JahUX/tPaa1MYoOPuJIv1cMpPDiraNvbjrMmVAsfo+EcYhuJY6PSWwvMhTgwleHAvc/YHgBvu+aE
tN8S8htKOSL1uhbMIc1eKqrBs/UIvgdBcwao+d0KRbelVHjQEYwb7ztCAEexqUKe+UDvqOm5LsaO
kO9kqCOId/K9zYW9dEE0Vveoot78LRv+qcorn2DK+q5dAcVN0nkdtglZ5wHQ0P/mWG1zzxZli8qq
Nk7XX7cIWeujFZn37O1crGM0XqW2ZK4j9GrAVZtiw0LC/w5tRUKVYysmLuWeNg5LQdLrKVwdphXl
zR7GFsdvwnlYdkhSPdqJZ3f7ce6YmCKu8X+XwlCUlpKnqhdjMAP1GyxczWbjz57J+8UO8ZUjik/b
CYymDwA+WHYSvHcrD9NqY4bDQlhU3aJRBrx4cHVnMi5Aj5JnFvTiUk4apGBDFrqufAOcPuiPEkTo
mxqyWorELI+Xje6ybfl8n5Mt+mrYLgaQTpqPEskpF28pSaBXRdl2LwOXfLuSw2nIXFn7b2Y18K5e
q76dyOUhcJ8KB9bw1zB7kKhSBAXN9MDYZvvjDyAaB/mv83C1/Lxm3PPuSL7KOcnRiCAPw6whFSWO
tGIYUXbEorkRf5xgyaFdqwPcK8l+lAtHcJoNUMMpYVS0IgNBF7yjl6JNkUnRcfugdDtSmdhWe2oA
F3wjJPy/NSrR6Wk4xMa1XYyxK7uoC+ttup/XvO9d3IKQFulFopFEZDbSi1XoiATe/Zy4RDKXSBrF
D2JA9yjucrBqTpPZGIz0DMneA316WIweA3Y1v/GNuFoZdPQIWI5sNdT0rNjPcq/N4EN+TJTyOQrR
SG7llZZLIHwDqEHmcXX2V7TWd/by5tPNjnhWt0bg5CkVnPmObNWvHBD8gk50hv6e29msjdbqin2x
Nw85hGurRJBqwR4viE1yMgYA9C6SCmwv1gBpvjcbjtIC4MMFA2IfCb/4L+pu080VBDSdDlFF65UL
k96syHF8XiUrP/j3xMGrKSZj0yLSJDSN3a/e1J6zo7NtA7Y+XfhLlej8HcEJHlW7h0oR5YjrOozc
yQtqdQTUeXE/xRmDfVoP/w/ABqeCvFCXCz8+byxpjBFCKEDw0unzLrynleByHdD9QSBBnLJpofZT
/cpwSF3xIYmbpSXcuNxCmiLGHl0r9tqJoDpzJgigxnygnkazWvp2YvhFtnJRVUGif9Q5mtpICms4
X7jQsYFFe3U+hjlD/Vt3iN3by5XXzWg1VF/Og2Nl2YPE6VOBPxDiZ3CE77IBJI4Nc1bJaxzUYqWd
JX9xZQMAbwFQKafJ4iiK4e7mQlcRqkt8bwEubAUDbCsfCK55K2wVRZgVAEwopaTJaEFwPZeUcsBt
xRiQW1OF+XD2lYNau5fu+PK3sKowsuWiZp4MqLfw74F2kN02iFDNLOmKYt8jrrMx/ygHeQWPX7by
jnqIV5A19kWN9YMFkJQQiIUYOhY0xkexNw2L9qkdh+/yeS89JMCeOzUEuJ+dnIrAE32IlxlJ4jpu
CRZS4VKVkvR+bSxrI2u/dwArc8RHnqQkSianP7rStGQS1jODZQ0UW7PWujq9DC2TT3rzDVULRpLK
nsG0sb6qNkgzsuHPKS7Kwp9jwBodbjHHwQeF64/RNzV6C1Kqv7axo+I5/roHHc1Fyha4HDQLnxHS
mg3v4dn1LvJ4P0EHMDlXfFDcVkZR1fKALKBiPaao9h4pU7QiAncCt6VRn9YqDgpJQ31opPnmCqPd
rgue+zQWyqudP5cwxY+Ba6q1fEqyAsTLVoIfBKsZGQ+IF3YqIoc8pSrGuK/EbYQJSaQJXd/r4zbu
e6EhHPHssvpZeRzvE1qLmyOwitV4Euab+308nv6R6uB7VLzteA3Uq/UMup4Cqrky739Ym8Ffaq0k
kiGSIgcW7ohLI9f3p7LmXjfUnwdod6tM564ebEEFz2sthbmA9rVo3HXk5aDlRW//jPADER/5PKua
n3cpIp8QlkBLX17l/KdTChit7uqbMbxIpFMV8yRuUwi6rBVOc42qsF1J2VuDmVMQSnSDAoJ6gK8C
Mi5T/wH3DJDoA1Qt1O/yrGyVksVjbgUKgbKuoxG9Czn23l3RlZAmfRGh/kWlwiXAHwIAeotKVc+Q
1YsC1DhPY67E5/FPdjN3F9IQFwL2ehTvOsuur6aDMCWRCZvaBQsHuXt2NrX5yEHQsUFx1UZ6FBCH
1SQHhuPiBeh1GU4Z+5F06l+mPJoJ6VuM25mPWLOCaq9wVEf6wdO53gs/9ffSWl/K1EwxhJVt+XU7
Zyf5rE8iZuKNvU/zCCARXFVR2sutofqw16KlkKSsz8FTFubuXopu0M5JlWGMaz6Kwu7h7YKJQfTm
5d7WaomvlemQgSlrMVZYpQTHyWJPXmOah5+z9v37atmcREgSnP6J38Mpj6lU+Otjxo0s4dqdGRUv
0mqDz5+MD4CQYIGKCMz/5YuMqVrpfkeNzIwrds0+Csf89erRsXtaHw6dDcMrNB/uQgZkMkdRym3W
HSLUx915CVjMqY0U4C7NV6V0c5JtWFHktLigSBvfy/vVUsrCjIyJiOAbiNjHi3RpSwykjcuI4qvw
KKG1LLyya3kWZQvMb2jfv9TKRmbZVcM47zMCLExyM/TDsx6u7ZK0AyZrFKYJhTUSWgqVjXlRgwPv
+/Ys3o5fl9IHz2y41OAymbgme4Bx5npZ5TMtPNdRePNj7rg3lJy6ngIJnGo45BeNubUIOE9UC2Yv
c1cf9yDyrcxuqLamL8pNHUVjwIEMd4uoT7eoWVDjsOyPLJmZYYvDpy/RJfMJGIInGWdQAq0cqiB7
LY9Vpc6Wh07l8elZcbL5vjQkVjsxeRmZuYLKT9lj8q3ct8pg4OENEnp1EDJq/oHm4VlhQ7W8KND4
APFdxFiLDYxA9Oq+hutmIk38btRTtT+o5hpitrBoDgsju7vsGcz7POsUWeM2vekBygAqTLOfJraU
Ouy+IWvVicrfJP2ZOXAfQLckUws3uevXJ+s90uKLINuJ6pJFiXYk3SIi0EKDIPgMdxZRnL38Eo4W
C8yiTiVuBRunqz96BVmEIYer2wyng9Iw2bJuT+iJdxZHd2vqAIYStjjstb1TjNMLAfj/Cn04FyVm
IkANV/1D1x7TptQDPS8Y7MC80x1SNkVgLG8TrPZc7UIL9GrUJpl32dCbIsAZfAigWHLNiGCrcaqJ
RZXIOT6aEji9inmlxCgsLy5IzsyvCZCFMpbXbMGYAx6hXx4cJ/Kvk1zob0Y3wE+yTm+Z/KRlCNT1
BfK2pp4h8ZRdNbA3337kTU5b8G5fojvvC4ojMH1TY90gGy008lcbtgYW6sKeQqsAmoTm7/H93ce2
mBtE5tS73pl2FfSM7bNoui8JTVY4sVQtwnLndLPHKoLT7R9aOYI8Uni7EZspdiKeAj4j8C6c9n6Y
oTd7rAmGoOov3pksNR9QCv9M9m5qaqia+Loe8IQef5RPK2ic0nkEVvQUxcv5+Fq+Pi8bH/g2R8uR
9B0V4bJpo8MYXpuexF5Nnswcle8p9vgDUtHdD55CNmMUuUtZKa/hwL0+a78CICM1Zhjt3YtKA0/Y
PgGTA8hrZwO9Vwd5r8TqGruRlqVQFxofHwfwnBd4uFxUEVx93rynkwcEPAQ2/M6oxHDK5TI06H38
7ZlDzq/wZGKWFp8woiIeayr7SLx9tsDRpvqBFjDXVq7/cT9RHV4o2u9WSRSo7nFGMIXE3DDfkvyl
IDxHjrjQUfotagyqDn3Gc9EQzd2WBNbaPHSn1/mZ6tdHc81N6bwjzKZ8b/tNaQmFWwJs/ombvjLk
Ge7tSGrfv07JGrPz8NJYqBDYH75CgAIGqqgkNS72tMlMJ+vY6EPmlOtxlD8EUyPIQOgDKBgXo5TI
k8NIdYp3cF9ZwjsjsUtGlHlP+aduMuKBfP0SQ8nhYd7Kpf+ZufwSQExpHtKaY1P7j6oZaZ8dWDRY
xNzYeQkbNA+Fj0Qq0hQTp3s50QY2vL3rbMcHtx4LPOr1qIFLI9e19LrVGSbcr2d308Vqxs3EDv3m
pzP6uGQKg0j8a1e+jlQilD4ZSaacOcHUY6tWAYVEjgYmRZ0ZeGO53GiyHWDi26BLKiFyDxz4Npes
p17ZTLf93199IytB45zGMnmMLz7+Ygzt16nsaXniHvmBCm1qHgU4hs9Gg4pE3t6uNklMHHwhV4bt
hSoNMgyPlIopEpBIYzVISUTmz7mJd5F/LMjmCw1FbBep50xyaqa19IDriSc6e707RWrMgkyOH6Qt
aL5CqyGjpqSNl3AZptx/co8N8SLL/jB0kLRZjv01F5OQe+zj1xg70qsoO/SCatOUC0F6Acnq2puU
dzHKvpjwIiiFRLUKj3SNngGs/fnVZTj2jnBLMVtBektzZypxJRofBH6lYCidbrQx7bjVrBFrsnf6
3Nzm+t0SlxvklOjwF9zf6qNEgqACnyvdu7kQbuNuN8+W8tls9eqW/mTP8NGd0967ZKpvQYSoSxXH
CgyxMLspW5NDPqXefhImE6qgs7kyNmIK7d8SqbPFuo2dn9wzWJ2yDIisv2JaNmU0/GQqQkmcam+s
aN48MZPpCDSikZYh3MvijRnyL7PU82uwv8DToBuTPNz0n5SkHn5t0gF7HBdXPJYZ7oqYnD72e9Hs
kYBP/OuiZl/AQ2XFlgDviSAlR8rM/UUHhiALWaWFELLz66AWaPZlG4y/F1y8OUv0YKbfadpE5AdU
SYdqsS33nLtwgBtGVRnn86BmyYzsHIB2op5msTzr/pfvOCxNdE6qs8K2kSDtS17zKCb4313us1k8
X5tHjGuxgzraToC/RxiyedBjenqsQTqBFCZS+Dw4RE5Ctq/FSi3InFoQPTBnEh7IUnOODprgyUWn
W847JnHK9JzhxxSTXy9+u1aDMHSLvlFsWWWbz6CXoBKplB675DJ2zGlcMRpo06grI2hBFKo0/VlT
BKdZDlHMjGwshaepZppdqZy2JAgf35sMWG6fg3vDc5TpOkNPUfeTSaaLHdE7qM+gGmthL6oTTpq6
PQTsVt6qmA/QCI4fyvtHj05U7BJuYfbHvTUdGUaMgC0W9QS2Cus7lNntbY/BS4eNFLYw9CC4uf9S
E2rEM8CoFCY73MtpR1SuL0ozNgPoqlfd21f0zOy/Mr4TcKl9oatGdwfUDpahacQhxan9Z9VadOR7
E6C5m5V/cAQlDg6Iq1O5nZDhGMlD+YWm6HBLkaY/osU4WwlzHK/hTMgi/YAl5qHmpoZwqk8FAuag
eHbTD5s4m5wtnvw2bN/Df93GdKTE+y9owIsXsxTBipz+hSkL2l+3rpBlPmOyazbzzfu/jfDBV9EO
PLMJHrisPGT84yf9kfq3fj2dkqSm8w/vlzyFYgqRIPH9x+CcyXU3Aud7v8t8LB9aId+bhHxhuH5K
4xqMNCycqXgxzkcRhkkQMkSvM33dj2nbusFVrCJUR9Q0g9R5ebi/O/URZnxv2iq3NWLlhpK4gfk+
9imLNPYB0DaugPk7ygjx+3K2kMDpvGyKfAa0d33WDqJuvYFwdwuwvRXEOvNdO35c2lbHxBQTRYei
tXz7kRtcNS9JvkZFT0Ut134r5Bdbd2uVHWRtbw9iUp1KPcPvjBzS9e9H1YVVVqlVEAsvhHGoqSOM
g6msCqqEDvGOtI4iNnPR7YlPPylBJdUlHO2dA8TEVDZXZyQtebXt4LpULpbxYDipE4a2XMWJH5P8
Ca//zvDpgjM0mm9s5LlXJ/RP7PvPbbxJoVrf3/DBhEmCoAOGQAmZdf2sXXxGTEoSp5K1sNXBqi+z
qmNpdbPe+AjLrhwUFIktowTqb+FNpkdD650uZ09NU7yC5oxfP+vLMND7t4Nsn42hJcIURm4vMS0c
y7CrUdanpeI7Oy6oUD5VUhD1HPQ9Ecwk5x/ufYp8ZKV3hDQF98uZIN9JVATaSCCwzS18Ff+oFErz
4HVwNWFtCFXrOhviuaJNGBqtAq10OWAGVl29Irj/TnBZqJ9gYtbmUDkbeM2p2fvlVix6eNwdaCQ0
2gtipKgrCWjrJMlmBhS1cL9ckkg9zWAxdFNRoNDL2VlpT8kQh9msBPniyDHvElfdhaecPI3r1Nj9
xwnzgfF5ZJNh16YcY0t56bKODkLbhGS3txNAoM07gqlztjXuJ0gH+MfPjKqjZk/1PtDWe7m27uuu
2tBjcDwsBvOjaEDPnbqWxx721HEu3gexZCt3NpUeYeV7qKki0U6/5/vUGQXCpwqazSQLoynxD45D
jT+1DRsCUObX+8geS68QZ/U1KGQ7RfFuT7gVURhWZTXquoF/6STwtGKtQdkOH+0By4HPqLKswgPo
72g5TTuQU8uiojfTkweRk9YOUqz/Zj/C2FOsiakwNE8XEjNHKKh0w0powOrWQUjDdGTgBjsmkWnG
ieF9UIajJQoKLPuzA7SwjESj/o7OKoo2qHqF1ieJ8rMaPOOz1LtTTbIatnWEoq9s8GIrGOdKGDVE
DneBfIDl8mxVFU9wfzlqGg0ckm5bpXRuNUn/sZ/Gcu9sCXxynxtWfiB67eQWD/0EMuzH7UDH8IS6
f9TQDNxsGCMDCqlhXoyRi5GFM6y93TcD13Cq0Wek1iD5F/07DF6PCealnQQREc/9tyC5eG5bM7TS
pp1pbiaOLyIb9XFqD7IBSW19/MSXqkyNYPOTZGbvV2KMPa5Y4pVayjZ56Yxv/OUwc1d1ql1aE+Et
2WRPIlm1dRkj6Oq4eVcWnubVkWEqmZRl6QCAAfD2b0mwfHwpAhpF6orqYRtUvWFfVlhKj2mxwyxT
nzi56JJn0EehyCsockqn5TyE34L6/CQe3VVhmsVDonV+IYmCA9WcqbnIAWgQjqUsmdI7b3PYP8xw
cvePkxzm8BYamoOoOiQpfBeOk7CtuE3FDvAd/pZK4ORSZmrEoR4MxKR3ijK36liir15i8EwwumRU
nOSkOGL5K/yTrXGeabrmHGDLu3f/2HTznL2d8HhhnnhHCpC2x3+OAO/oPKqwDl+9BGBckwo1Sx1o
bp25ENuJT201Lf8H90+6NnzZw8mbEyP3A0nWT93cZ24H0IO2iyyZkoQhA3JkOcEjuEnAbL3iYwaI
6/lYp3rtsQUNLByPpDivJ1g6Mm/WnqZqax/UO/PLOTpJLz6SrcZM9fLD7pQ+/AAY0zoE9y00wg7e
km2Ky/C+I6uMd0gsHUTgIhChSysgH3Gl2Eh6GR0Qq8XKC8geJI/9aaSVDXun4oSHzQMZtjckZQtb
e7+kKI2nv/KUMkU0YKvQN7bqrdyvt0WfnIXrzY1IQhc54EJrUR80sSlG+kYbQ+8YY/uja/8PaMKn
JiBya7atsl7ZNidyYW8Cr2oUzcj1AmXD71eGhItHVkC9QFwar7iyzdHuLApgxPYA6WYVqxJ9SDPo
zgxyp8HVcY01jRI6pf9Yz6y7k1+c3qf51uTotEhfR/MdQjvU6vJoDkDCBbOHK/kHKckAKkPIUUtk
VnuyzWaIgCB4YKFCiifW8V0JvhKsQ1ul5xyN+jMcOnt6lCQRRXgT6xH6by+zbWbp9JeER6pdPJXF
kk/0pcPpuVJT/BKwcUOi/8OZUgN2EBFABDBC12PtwZqG8qGGj1q+4HusPwUAbIueM6cPknYpKXkl
FQehFQSnidsk0QCybyGuBxWFRC5LtvPMRUVcYC3Ahhc+uJgYnvoh5TdNGwMAAz407aFf9LlKXCrg
2cyHF+npzkqA6G8NdW6shZHx0fb0h0OXJujk3ZVD+sbECyRCoiRq8yOmu6V560cHiJspIj/p6FnE
aG+s+MFMWgmrWnWazm+AcoIjxBPaHTev27/wHkBjnwRx621OYIkhN5U/srH6CgnDF7udn/SCKUUg
22ywQ7kM8wz5QY2CIQ18nI/W/PU4qi42StGoB26dXyi1ArYGc6dnXoFaTd8a9mlMoLg77ogvYAkj
8QuuX2mKSnsG3Di4X0DB7jvdqIyLIbbZom4+Ld71FWWuDLqlGkxukqU+POM9DTVBztnqVLzlMaEc
0sRxadkgR8J2KtpW4cd3D+ovQtoGN6zWso6Gh2VU54QhA19mRKqtQaRt/FtiIf2D2acYlhDvZ/Xv
8j6Ynr2IpN0+X4ugVvNlyOisIyTtdj6Zqd0lEm+qGZIRdScwyRQgVLHBOVdLLMqhuR/QHL3hx27Z
dXhOyUadI6cbTrHqaXJ7hDP/pKsHs57fp6KuuwNvVpKAc+XHBiMtZAs8A4aV6XfXsbvi6qRyW0/w
Wd3NFnKf1Ch3WVaHrr1vJyiESVlB1NLGscq0GJE2FxioYxnBJrpohYiSH6qiDCbiRRhKBbhf3Uos
pphgIX8s+8t6aDKiOuvftIo4rGmSCv2zRMI1k5Bk4RiXFl5bT/6O3bty0SqQwBVk61YxnFQXnk1x
Yv/Xfhs7r5f5xG9MfvBx8xjvOkK7IjzuaJNWdYvpuysWHllBem3FYHcgK8QsYL+a75MGXrA9AsUC
XXEm7wkOiBkyE2VJF7lKDOiOwUYaC1pKIwb13VD1It7sBSnPElaPU17rSKhtuZPC1OF5bqg1qFSq
QKc63AscU1HvS8HgtfhY9I1RgurH5s29plEhrhATC+oknx2BFf722gVUugV3I6CU/pay7vazreQR
3qDylEzy4fXVgAgYESjvcNHrUr8zmrev5Jl9u6lcqpctUfWNQN33EHvEZCuyMlODPF4CNzT8N2Ht
IUIG+gDp/oSOX1SRcM4LEREzfVup0jEeXsz/pvCO4dnya6fzHGVcHsgciyfvy16ycovruOknAkpT
SZWsYcA9P373Sh2gOVhlldwumuo5Bm13Q7zIpJKtkBf88OBWiGdczTYe141b5EMVp4A1+KW5mjg2
KuKO1iSPGCx1iB/SwoMRrRgPE2QmXyy/fnZu7QSmhwFUeTFCVf56Xq4LVqBIufttIrlRcrVbRl2Y
VG8vA7VVHlM7lj7h0zZMdrBXGHnZu6/fnxXNa5NwpJPUDxloSgUm95QW4cyTgJFlI0B6ljWAsAO0
EBuRr1qR+/DB9Flxhx5dWNSP442jmx1tDzcJyf7l/3GkrmrAbnnlz13Xcqy95xUzP5eRhUOaUjGG
NawK1HHo9HF2VAuvEoq1vaZ01vW1jtr4ood1FbPxT7uaWeetKHP8cEZBsuS+lFMPKQFRraN0yfIZ
c45RGXw7ahdnP5XmTqd8nBIoDenu2HUflukjX232Foo24iH7/Q6syj7JG/ntxntg1LGhpt3m2J6k
oje69U1iuljeHqd+NMpJMRVXCJb2mEHiY/tCDwzVurm/5BVGFKLV9WXR8PvmdxNiAhUF109mG9VU
OSu11ASgP0eTlhOw4bYYM4m0pi5Y3cfYwTUIl/cnROVRqgffr6b3XHwmBKDwXXOzuP53OsjPtOBt
qTMFHYaidFGguehGh/fE0nkDTxLaeSh0wY9A/ghqWMzyJ34VXAhXDE1DHksk9d5zbYSNkfJ0RF6B
qHkhIxJGmkcfngteqiLy+dRzU9J4Kjc3qpgsGSEIzqmYaMjikwCdS/oS/5bC9ufS0DLsfbJKszDO
tpNqaW0izYZdb4MyXMwabEcU122fETLI/iY/7K/PtTEKuead9rt2u+DwxKaQ06f/zvGbSwGRhD7v
xFGKycM0O42dZdc00LDBkLtiSkg8DV6x0P+zlbkE+yKbJWCESeMWU/wLmVoRsk0haBfOa8n81P7q
wzjEQjhuRWRCKEFPnXSi23ImXmnzmUQ2nDdBMilnZhrxRdKMG0V6R1Gh54paRlwVV8/tZum4a8gH
q72hzR18JhVivQI8SpzAYbmFrnXwpqMDUQBDRAgUCkjetcsovaywuQfE57MHmAKynrkNC6slBzHd
R5lzZaLSaQl70R5v1wtrh06a8pU+oYFprJipBGKumX5CeV8nuDMXIFZSu4feSmD7WpIYzluT2Hq1
SlNVd2hrxeSXqBjJvjWm+5OGGkGJY2KuBV/GdsjSFGBe+B5tuw0ZhgyJQ+mLpxew1avsGgLZshxU
T3I8RZ4VRb2BON88NhvRW2wg8UdHbI8T/kx0drYd7lf6nyb6WU+m8SUdNLI1Mx9ZXKPIWmI8pEdL
Uv18/ss62gnIbsQ8Uioj4R7ohEra0bsRzPEuYOWfErvEypbELj1sq4qkPp/jxmDBEKYM7exFCzbN
iih1ey9aeo4tMkkfzyRvh0WFDV4fy1f6tvaUlh8/6z0fwFniwb3KZTIDkRM8OXScy+HRlejebWaa
a/uHuHZ9yQ1wxFdhzzJzaRbQ/N5LGeWiAE9F3D5SrdlqHBSi2V6f+hDStIzm/SvIBOU66J42ffkH
BYyEc3vdfMo2tCfNfMSXHuhs8EIWeRsv0dGJ+8GfEhJKl7Z3vxTT0oLkDgG/qbbflsiIbmU9m0aP
IV7HQ3fxYRvBlac3QaKvteTs7i8oGtVKjQFzN0VwdUzIDPmvm1chjn2tlgLiV9tqmIr7TMCYVXyp
aU3CIKGOa0JupJbmLtyhPqv9xst7X9ZbPW1izxk+F+vmdM2HIe3+XNzkqJcYkLlBEFNozAOMKkXQ
fWfzhcYGwFkxloEw7GLGgpWG2uUuURi8dD4JKbUJflyBHNcX8otUXRCVuhBY2DBkQETl1DlCx+aP
179ppMK7Ic5Frk9jHs12HKKdykURvGrUvQYUgwXgzFXXv9QAlFozWZ7BNUlQ/XpQhyBynMhIAIua
8gQNu2lkC+DSW11qGjgdsko9nD2nL13MV21H11qSF8S8T8tvgNUDnCazGTsz/GsVb63re1gJWr1X
rOu92b+zQLKfQ9KEN+0FeHtzYOQTPEdB/pDDiGLVBYfsUF1C4YzsAVixJrYeY2p4/g6NOT1+r8Pb
YertT9cCIkxkGRHLuHdYAGdqlri+UKoJPOPZ3vtKYmYLdxWpR37zKWfGeZrrHDZQLlNnNRSIMsLE
ciCH5zu1Q7+ZTFhn9488D/xSUUktD/3FfkeoW0PRUi/n3a3TWA2d9z5C3t5h48J7cehIL5E43ols
N6g+XxtF93gqOF6b8whmbP9dygKGSbkK0+W89Xv5AmUeHOD3fbI5u55UMh16idtHFMoP1wHhc1Os
nEa1nZX2N5pExUJe5iuvrWflen0I4hc08oJCv2loSk126nFnWyMZxMLxa1LGdrwjZjphxAlqAr5i
sZ5+R5A6dSFpRQjl8eKUZEkAU92pBKknnIQcn57vG3RLO8Q6k7O96l4sXq/q02Zs1NRWB4g8vwRf
2VCDV8b1n9fly52+ilrFSobxf0THDsOg13rC5QGmB8guyJ6ZR0CTVt1nQFVeXT/yS9QUovN70XrC
67/FgOdslK2d2H4VDNu7/qJzTtHVUb0p1IxKdRDVta+P/0yf1aGNwdoKOjUWMEE9AyJiPLDXBgib
DNXOW+BhB8rj6AdYs1iC2shwNJSkqG3UxB4EKmqkb/usaUv4+60f+m7Ss9XzeUZCBdCR6leL/mS7
dboYbYKGRCTe8DTOdpsaSId47+7iQRtPVREiUhGo3MA+ei/i99OrmNA5cEL7PG44tWtDr5gR2G8P
UOQweQ2NWQo2IgEU/CT+iC2TS+lFi+pTThM5t9Xt09a89hKIoSBHT+hQcbVIjlI9V8kErjURaPTS
SHH0bR4BRKktABxxrEhGzHcRAPeQOr6ZU7VE5c2cfNNsE6lV6kSm4iqQ5XxxrMHko47xefczQUGy
SrZsgLt4P6A3DE8r7bwBzE8dg0LU2m5L7hCPvj3qo2vFUrXmUeK1RbQGgwcT9D+JNrFq+mL5+tRF
jhH1FTUauyEQw2XH61elY+BZXkFpMmVIZPTbcu2LBhrWc4Xv6A/wEOzDiO9F4Hd80n+NZoCG16Lo
hXX4LuQa9gdvzHf8IZxwX2SO8AtWRq+B3SCsyJG65iS11g6n0cG4FLgA+LCggTFXRXsx81l6K20L
EXU3QGyENv8WKdvNAI3gAi4zb9nLAVyR3SOnw83pLXPG1coQFspdVocEDHUmJOvOIW5vMJriJctq
0vRNXGbh5eJ4kKUl4prP9rfgM9ovA1jl2zkiMX3O4r2Ws/6w31jaQTQQoO7lxVXmletHWnsu0Kyd
MgIOqrNJKKUOcWMqUyaZ7S72gPRka6sorBeXuJ4W/ocf+cXDcOVjnzYR7euLqivU5A1z/TlEaGX2
og71xERgcIYvStnvj2PnHrDsAeDW9Bm4sJ06gSSMWGor8tNIIHiRoQsILHluInJunM0WFiGwgfnH
ICQWfzv9BSb/ND/xBbvHw7H/ZquAFqboBHXKL0Lb6OZRJmhf4smlMNuRdwp8ZXMvhI8LJbB4peaK
L+s1dKT4P3c1+cmroYOxwdj1FmbyZnh4tuolRsRM0ELugVOcqc9kcYZVGWqsVI/08+Rs3ynvN5To
PZ7p9N5XiaLwDYnMYVXjbC8MmXWJ05ntkUKlRd4G6X3ligAdy0R0rhV9rnF0qdOhseI/GJExIrtL
NbH3ED4jpbW+d3ogIr38EO45411/cfDOlzHum+79vTtC087BXf4Wfn5KgBxncVlVpUm8TwCPczJQ
Dt+Ol8ksIDQTChQSMUNfD2APiAAg+ltXgi+DYu6Ieb/Y1/sPx006OYar43f9eOhxD2v/nkLsjsYX
2itfNfIc4gAqN350xuCNnue/GbR5u+79TJEZ6k77Z4jAUiJj7vBZXurwI/tIxqq+fnTNXz8NfBhy
Bv4LGRY5ZJbAUFri21jrb/iKQez3KmYSm6sbJbabidIl9eJ5SIe4gqNX0mKliWyqvz/WYUhLApLB
aVF34PGnMLOg2T38P0ylP2CUxWFfLZseVXebDQFVxM2z8e/zxJmQ5ZNgMJ+pnRIALO9D7jPBxDgJ
I0Zpv7BH81naS1dnHdH7FChFlIFS/V26z83lZiiYSJD0gFNXfxWdUsEVG/trDjDybdTJhx8cbhL1
/6hO5qSAb03MBEf4a3Q96Jepn2ZpFB8M85ntJhqcGJsRNJ3gAdfGw5TbRh2qkxIHRhlLN0yemGb2
CZudaPyoGQSrvlKxca/nn8k8KU0uWl1bwXkP4WMy1XaKFlNDVFTCoADCtaHLuhI+XGXZY6Pf3l68
cRHqqle0CWi8ssadGyhlL2nxkYvxhFTebE7dQfsfY6Uyc17h4q/93AJMraslUurW4LpZWPzekNqh
1biOnxpv0GHpoOc20t/E/Uj74dS55RlgxWCSj67EqZwd+7s3EgSc3j7ryA5bhuAF0Q+KJauzwBZU
DriiXiZfXh3A6ZWxNWD0/KMkr2Heln5uh0JyNEmrKYDK62schIjUH00xfjTkTZzeFqP/xXaKoEfv
t/iSv7SuwaXiot7iRw2BqLtZ37nFhj6Gb4tHImkHI8bk/Q4lmIpb8dn3KWqOGJHCAhPS6kqKRsbG
+tADEJ89SYSluMjzHbvMWUF2UBCINdYiAO7IERxaeTU4P3loN8pWfzB3Zp3up8EvBdmy5q2xUQnB
zujOeS0O5rx2R1sK9H6tJ4B3UM1gR6gHgDjcJYRgW4uyNMu560dxDGv0sKEvGnP4cnHFVZ9hwRod
r1MgB03yCXoHCl8tWtdx1y1mV2srrPsmFD1myWsH526Cdx5ItDvSdS3W49iQotEkzrGhddRP7EF3
yOucEWY5K2IpTIt9sYG6n42U4Fm0/D+kqzixTTgKV3FdGq9pKf+CfJI4D1z1hZlU1wJH3k3Im9nc
Q9nUCOXrsf/3laOjgfzBE02jKyTDiJ9c0wO8XVwPBtsddMXBKIMrDmehJwZUOwT7azX8mL1pQa6+
MPAsyxIkRd/1Nf7vM9XTMFwEAe2StKGvg3kePaPR5FF+VAJBWGpLb3kfkAp7z50odW+mRx6tW32q
j1x+QkcQvALgK93jlx7ES6ZStNA9/ENnhV9qM3SHgGuAGijWy4ur4tOAuLE4J2QpEt6woOVPc+pv
CaR/D+Srn1FeFKInM4ftUYNZA3pS5+3nhBpK+JseyLcEARmDPgA5lpExKCknNAR6VCyG0YMb+ZHz
MFA9W+GGe0XdRsJCTgwCA+JO+r8EfeNKbJlSuJh1vwQG5Ov2r5PzG0Sh2zQ7yui+jgFxdQkGfEPt
EvV3P48uMvKmOMHC5M6leQL2Rn/Qvl8+ebYMumn1AMJYzxU/5XrNpfyiiPlXBvoQxoEvEXHUBmLe
0/xqHIOw08qBAKuM+x1zhdYc3fSah2EIZ/rXnPq4Pb68h0W6O92xNf1kQ+qCDjpt+xAPJhKjtTBS
/z5mZ0dTmpuRoEx0Fqt9PoJ2JrHdDnr3gEheEcasaU3BJ47NCExhVHZOlwuShcwK6actpMO41RtW
d3/vq/rK61jgB9De8jUKt8b6wCqWGqgfB9Nd0MmboRyDkO5uwhwI7itOPAz9d33dVI3/fIL8poPd
CT1zq/04SWqbQkkjTmtI+sQhw0aXq/Y+tBSFQ6nbgodjqS0uWi1mZ3b4tYVReShv+zC3nuxcER86
bqqL7tulSreZ0Bk/9RcTzVnYC9L1YLIbVrOQbpQ0tHlk2MN10fMYHdOmroXAJQTGLHQyRmUZyHda
RkCcZN57fzTu1l8AYZS1eUBG4Y2erEQMSeCvTtIdDP4uLD6W30GhuZkr8vOy3vlbflh1G30bOomG
DNjNRgcgo3sHrHSsvhNy/CslI01K0plh+kjo07Mhfa5Y4kcB7/rzXmKhIeB+eEFKTD1zReR7P3vf
0Ad5k65MoGLePm+o8XtUHXeyd4GNoxhGEP0dXUd0QU9xB2+vYfOqRmJgjdFI5AF8CAjt2HJ2sY7u
1D095gKLFFYj9nIhc3C1WVIrfYFmhmZvpOW7YoYj0Lh9358L7A8MImObyNY9Ctg6K4KAUrcKz8ti
I/hLRMVBcXK5oBVpfhZZJZ8XMcQ1vEGak/jciBVUY9hBNW6sW21ryWOromSBMA0tdNNt94O/dUXl
9vBeGCJoB6+jyzn73R8PpHixcrLY8omxCiNdvH2+M4Oo09iEnu6QooNGx+MtJZ2+11oLXhOYU/Gr
HzfMbIe5ghymjQ8rAa2GuXfFitNI3ys6IokBiRAv4BcOUTUVdHFmSfTVPUWnSNIKnTV6orIUxbUU
wf2bHkQTBAdDLDVe4+W+Nky4oFByhy6ptccmeWt+jGphqex5U0mpq4lINCgBSm9ntcKeFVfsV5Kl
sHi9cZa+zBl5hAwVhQQOGygwJtZ3XbZnWLqPPDWpEoZv755E8YKwydjMAs5PVhtNlTnPCyzx4gmt
yFnvNwge9dFof07RJUTv6xjmF+prsGmYbTRE4E+eAW7UPIIKJM+SkWvruyBJZscKTBReLupD7gjW
/19GvI+mP61aEu204bspwQw9Pj/hK0z7cFJzza29Ds4BaaAajkiXc22Lgx/c8ekKMuVGyo/5wPK4
+fzBwEkIaXWLCQX9RKONSKHUYZkhbLV4lr58yGAeZzOiNVemLTWvRa6neZQpIbVRR6lnAWwi+FgE
UWJJQS3VVNR+N6M2F6KwBVcFHzBavYIJ3tNM3kJ2flmJPD6G1a8lNEu5am+XPrC3N2kCd7RoLB2C
5xNOQxhnUjhGWu9DpDkgjSCCRXMQk/GIfJaYsLJCcPz0AiIHh2olQLIF9mCyv3Qf2TUttYRpBEcX
d2r7duxoJ6X6u3fMlymE0mNAwEiFia6aEnUJrVaEYfM8m3kC5rOdZMYGHMU/gw01tFRxDmxQ9rNU
3rgTiQe+Ywca96NWgG+ZxeCVVujgUSUiaknSfqOyKXgFnKzhwuia9lDGOqtO/OJhwJ16+uzh/0mW
j+5SCcHAk+K+dKk0u5awwB9murQyjeI5AMifegYwUQi5yea9BbpZ6dH5dmJgwubUTs5qgtRqXjUl
vdVuQCdHgc+hNxVb5B3m/RlUretOb4chEpv/oEmIh1tDJGBWYKAYVEgVfUQ2BBWns1PsCGEPm3cZ
z6RDL/bN/m+lhI23b+tauvjb3lGZWAxeGVroLNJTfCa+hyOKv7EwJKlRSkiI04CVwDIj5PuCOmjf
3T+/DT8xNQRL9EuuUuTGMoaeDxENosg60iRNvQkneshEOmRJMPq6ATk+WtPd/A0RK4LNMLWAUadG
3BtHgmFh+zIo8w/OCfkfpjXC6ZSXjKd3d01obfbQaXnqytU4ZQITmatLH++cWxUhL+jJe5dxn0LG
0uNuJKiwfXD3Sulemtu5MaXbvNl2YVgCM/wsSBbSKRo2oYs+SnxmgV0X81cd+alNOha86jD29pr8
Dut0o4DCpdrDyjaQb0QTD2T6MS9LoHizMQ/d1V+dZu4D4ZQbS4XK4y92nK+RhmXhYCqRh4iCBU06
cRxHpUbANPkgaY8d0lbYnvYDv1HEW9mLZDz65+vAHtQbEhZqIP43gGRj+7MjiqnGaGDGA+4/VPJ/
qKCVt/fFw9SWnFnQqi9sEkIy2w9xVdZ5xge6GET5vaPJKM0mAosELWmSGfBVSHwGYrzFELQnzN0s
g152h+VRyfTSYGc0EWFQR6hF2uY/wATdlwXVEkLgNgfezu3R5AI8ybRHgCdD+kWclSn8inh9vYL4
wDO10WV3bSxXnADPFF1YpIYpOTz/ZH5xI7CCy6uwD797qRzM9ESW1hds50aFADT6RMHuBp6sD3Y9
5Ivlu+71bqH9RugW5/s/A8DWneedQZ3lsv+Oj5/oDCzQkhhZHek4RbbmL2eFMyOLyOQ7wASSv4+V
pd3acG3fE9cUKX9RFKRLhccZ0iZo+NLzpXhqNGR9kobdj4qW2q2MGpfnyEiHyTVLSR3thwz1v/Q+
2GuUwSV8coOPut86aLLzzY1NBi6+a/bNfPdz+fOeDCiBTrQNNEe+O7KncKah59rUAOIJjYHjMB7M
g0v3xUMGnGQ+P37RrMazdEihZPpFfo3t/wYQ+CsXwKwihEnItcB5i2GugfIrl5tie1UyvPOYQ0Fa
ovRhwk802I3mecJcqY7rsYM+7+1IG55iQqPmVx2wKGuBUR5X1TXVM7pCN20OkHZ8X8SmUYnF1PmP
00wK4kcLAip2b4Z0hbdUzDpqJ/dIGFkuUDYBtdenTdDrNhVwiwKioiU5MS+9T2kQQkEg9uUH83Uo
XFLUobGFNP+99B9PX2UHFxYghO/+4EjiK7TlpLbEl5BPBOD2ywVa7KFVkpPVdBm90TYf6lsrxcEN
Su3jZH9HfvzYgW+p5gGPfInBYj3/E3FBjyhU0R14+yBt2t7Em4mBh5TgAO/QCmyWfQ++oLpEpPY8
W2feMdThHgvxYSg67k36CFFthSfxCydEo3okRMmkDN4E6yM1EAeMSMEHVrbux6Sq9Ke0cVc8Kcdf
cmITNpMDsMEcqqS6LBSZX25n/kDiWzEAYdgUuRuf2z2BHVczwzP8hhTHo4d1ji3iRXCzx4uLiBJE
YAxDhoO0d8YR5LSDsbyF5seqJDSr30UWUCd/znnv+Vwx97UwWwBTZr5vq9WVOaFCU2iu4Y6o5Si4
7TGV5dIZRiMQIiAtfd1BMkU67uKd8UiN9WzfW3C3nuy7ZMP1kd+Ohh6S1hjFnsJ1dERck10FIOx7
0R0/5JI2/Z0pW7LPvEOPG7fcVeON3DSZk9sEXTyNR/bp2oex9JWxyFLgz0OVfVVynTGuJDDr/P9t
bB6XRK/QJPRt6NnsqR7RHscsdAUw/ox1/q8Lhh0ooaXRkLp4AKUsK/zIvCRdSAk4ex0L0p87uVTE
Id37yuIE8ZVpGbdpT3lhFlUGogX37Fq0V64OWXsQYXAlcaBc8MTksnFdAKQnN58xrLYPlyWMl6Fe
HO3l71ZSva0ZGre25aTcDxuCmdV0t4v5qe8cvpaNLmjMpr8JAEOgRzvR3LXUGvC5sknpFKjj5fXF
XLaLRRU8nqCCAEGsMs+F90po9dMw1ngcNfOe1GOy+rKVroocgL/XcMCYBwESJhvTTAeY3FRBdq2z
wdzawztqxx4W1qkXAX6E0zh3isOmJG12TMTOnsR9rN8H8CSbrV8z/c31R60XTNDyCb84Q3YStCIL
v2/u9o64TcRLtb48NhoNVa1e0AnU9nFEfAosbPCj8KQXu0srMBmIybr9sisRyUOzZvc1/YZdo7W5
+g5f5av+77GfYQ3FbTy7Lg0jjlZZOAOvkz/fiLKExUyy5p2lq7W0ZrkQsFc4aK+uOayARMSO5DL2
7IcvnKQWbShAnYUWwQGOhrH4t9VQBQeferi9tPaZDUkdtxocdKL1aJtYvH56334pD9bHOv/+crbg
H3GLaxx/sAMwEXADzRCFnQF428sYqRnpRB5o3S3DK52/UKs/aiE55DDOlHlnjmsDqKdHFWE5yikN
RRAII6aKPEZuiy9ViBBkbkhKiXpvJfLcv0XyZmiw0womOqbbhdbRugVB9oF3YG01lo1LxbPD1Rf4
OJK9m0e+rFx/dW9U28lev1iH27zH9teMxrBi0n860gq05ALWCP4HFY0eU4O28P4Ytx+Wpcrwzjm7
ellhpYn1sBtca48tK8yOJX/lKYrExHSi+cUqypYy82/ntQGI5Ay9Me5E2TD9F0e4vG/byuSMjNOX
5db305grwqEu56+dr+Z7tcW6iBaUSEmtwdycG/NVAUwIk/5JQn/fELhl3emb967KuXPWFMHBwLOQ
Qs1UxSK2CmNshch4QF8wH+gvnIG3BrkkO/v2MqOPnID3wVjPtswWRPikw0qy5+4wgHi+nK2UH24N
4gqOXggT55KpHOqX4E+bePqN/HXBv9MTbjJsKTQ38PZ/Ft3GqagYMJ1vvEe4TpAfiBv95SGAIKYz
wCQMvB/sGINsae0O4a5HLsK/ZVDVB3hRp8N607mBWLW1zPoOmtKwG8INd6vUGZp/eMsfsW/jJbEr
SrxaiW5DR34HJNrJKXgMy+rRIfDA7WsK17fE7erkaNfNQm/mytNtDeFe5yrvjU8Zw7eRefDSKlG0
8kr7xmu8s6k4bvkdl6zKZlmK76wykmdEelzscBN7W8JJgejnNVOyIkPV53q968ZlAEB0RkcdgA26
ITMmwqqYACp/R/4TL6/egu/FZFenbkgylrRmT6y4BG5WD+PzS05Ijp95iXJ9IpIaLEQbihRd5QjB
60E5dxR1zxGMkf57jV/Vd1aoynjAsX03UmOCQymFTBKx17xYfvYKh/jPPhCxlpFPcXd3pysmYju2
JIIXtEgB+CvHER6YycYaT/uUkJz1bHVu6V/PhwIlePjjELvEgqoqHNZBMnXrH6D1Y0fJO40JJ/o6
+tRFsMcCgya9A+6UdQQnO0yUo4L0Y9nZrkpXtKLDWbWsDz5nC96LUjJHHr7Xicv50CX5SuzzHR5+
4EiJineq6YxuHvWgVizudndNoU1aa+AH0EDF0QSDPiWCWmf+JskteyJs/pgeFO/2amuTm/GtJV3s
q450xZl2qvPFLzvQHJe6x5T1dyo8sxdrVosYFiukEilf51DSn4TLmmMyYiFlOWryBC3J0KRu+5j2
/VsTTvvbrILeKXPlMqSnAaDeOVk4UuRjNybeBHkZExuVFR4VyWx0v/PgfZgz+WcHwf+IQ3oSY82F
uEg2aw1z7LlU7TlQQBHtUoezJcouAIKHl3IyzsZ7yZdaR502z/lSAW2jf9F8dW58i8dCTWGH6axv
NivlZ4Mfe+7rZfX/s1AcJuYYtMIQn/Xaf0La3S9LBCr7XOpMG8PXFKZFRZd30EjDiJXThAIMNrOe
awsgQ9cSexSAad4DwdWYMg98PMieux31LseZKRFBzbKJ7kJUSnosmLPj+PYobCQJioU0xF/Ikq1Q
6xE5Q9cfb3UiHjfT0p0RcoY/oRWmBl9v2Rg1Qj4GgTeiWInPtXUV5q7PAwj/vJ8zQaO81BBIzp01
ue73SHbJuI4xTgKgw66e6cXAnJzzR/9fGWwuHP32GA41Dj+G5ETMsWnoHCW+8WQunT9qnoSaitLG
aadgWdwbOZUMY+zGkA4SBehOyQxVeJqjGvwJ7EMRiyalnCBTLsV0FBt6kCCjml9VptB8upSLzClD
j32MPfQMLe549Emj4uLEHODMa7lYO/pO4B0eEGJ2rQzFh0rWttjhuSiWHnwMJen+qfhHHYP6BS4g
08+HlfbpM3Qy1jK8LZLOWDTWhowqg9Qwi8GYWJb+3BiVYe+NkBC4cJMqcsEF07rAk80fFJcaekzO
uHG9rk8KYaItr2d1NHLSee62xQ4u7kcxJcL9WdztGCPU01NaAYa9Kqv1IWZHHYvm4wPBEPzlgF/l
gV/juWXndXK/egojDVE+tinndBI/kme4KjFQFbF/OvqCPbxrPFYPwI4NJ2ixnGwvUVWdA3l9bAmE
RlZyY9jKgKtnvCFShlE50mZ73RrnVgISZ0PkFIu32ymvsPFhXcA8o3uy9unqM1NIXRn+TZ5xPgLz
1fFI+lf5rXxOlEQG432YucG0uodGhorGS9FTu11ARd+iMLodgI5FZRTXAyw+9enQoSA+Ff2VMBXy
iBuAqNn/XHRSWgioHU90wiJwwojCSkFlDDwrfSLlIdxrwlvWJNycwXKQQJx9BXxOSKK7hAxCowER
jJ1U5kyOJQV31ph4Myum9l1hwQ8EDP3xCqSZtodXNZI8xvNhBHMiIwTw6WNwqynw7Cb3NXnqQCL9
3pyy4IwqRWcl8CZgbw3udFqXnrpg7KLbvO3Wcz+hOcnMtUoqxlReqlFSAkt/7KGg05irM6RxWpAy
9sTuwWM/XNZZiI2KUe7RIWmUixbWnBKefzJoloyO1/q+Iul5PofebeDHpqFC7vcBhEu6rlNwYvgK
uymOKRhnTeuwMd9aBb/sYhEBs0d6HkrFFD6nh49um6cjnuUB+iEOVAy8KAr9hx23Omp5zHADV582
ZdGIU7YhcYOYSTgX2MaQKK+u7hzbWZXnazpjp/Xb7GHo09GLh8Ji+ncHZR3RGxL/kzAyPmojcdLP
Fk5qAPuz8GhviSp2ssXQD1skANvjvmi/8Exm0xGU4OapXdr5m+xYeeYJAWSX8G9ux2NWkZFaZDdQ
DbpviMFfTMCqJYQfHOytN9dt5/stOlbCkQrb7s1wz9SQcM5bmDFHee9tbNT1wc/3lCDWG5RN1Ypm
dTFZRN2tUZjQ9sIDNnOttHlO+StooUd2DyYdZgPbA/unl7FZ4bnwKVZRDltSAvXOo4eViAdpRXyC
jwDE3HIciBkvk5QrYLLiszRHkReUEqPrPk+BSh+3PLgr436mgMlKi7+gnrSAyrkzAy8yHy/2IYue
0+cLholJ2dQDf9D4hgd3W+Kiac6f35CqrK3yoWdjb6N291Zxz1i+93jiZIyn6CaCIECoCKG3zeQe
Pq/CU15F3k83p5Mq4dwiNpPqp0C5qKracRIUlUUortMoHhRdl7NE02VVticw0e/MW3JYR7RW/GRK
/PjEbLbIlKTV1s2NU0p3KhTwwRTkYGPt4URlKMddA74m3bzwgeSAd5OLf03KA9tEQxl3tD5wK1ii
l1mO6PfHllZ2/pvvB8Fuo5iXspVneqFANMFMI4ncD/+5+ViCeBs2KFN1Q8GlHhAVje8qGhsb6ITj
B6+muAUTqVsC2WPTJYEn0fQbf3nHxuacXf0toIYjxiET+I+So4/5b3CMO9ckVGI8Dn7l8WBzmVlh
b2tykcr8rLsVjsHMZctbP3AFyoPDw4eLaJczWK5/gO3Kx9KICMK1Oc43VbjQM7Fn/BheN7EBLNvD
2EAd1DvFgYwx0/WvHHDZgVO9wqzZsv64Myy8iP6lr3Hj/EctA3q4ln18ZoJLmpEXHEkVYDfR71YT
b6Llvh2jiueGR4qsg9lVX+sKHuV2CHyfnUu76g5YRQnQud/A+r3U41NTyani4PrMw7t+HQ3jnkw3
GXPrrSFtiAT84CUtHY7PfJO4L/je6yGe8f7rTUSykDkKGiOKQkSlS9wvvW96rGGGYTLzqtxH0z9U
Y5M2KIpxF0Mq6RDVzSdNp5gkb1Gt+/+Sqkv47xXOELzrZYojheIms+afDg0Om6JFgvmAf+B/K7w4
j6nlHp9uh0PQob6hbkEhO7/poEOATMbcknRukbl7SPQJvnD99cUVYtYgT1G/fXwYtzXbpMka55Jy
k+jPpbD4r+ZwlNBPwmpzaXxpQPkfauFWJwhmx8+KNFzzTvWgy5sFPymciw2qcvlYsvPbv0t9TE0s
cAqMQ8c7K2fa+tTbWnFyB6gR+9R5eNphUz6lPST0ftpI5C1+pSZimSuApcIClLVsq6Zd1YAx7bfO
NZ63ZEUjRgaQkJYHCr5Sw8Xdb6vFbvsUkBqMT9hp4EjF4kdQ/yraGLSbh0CdF+OeiWMPdlFPKdzV
jM3l6mCRFqzwpUdczXDch0FLub3CuRBTdAKPxOKdd5RSPVPXxnsaKWBnfQgX7pc0eW4PMOz3F0vt
UDX77qr42XFitqDxLWdahc4EOnVZ/mAYwfCxoQWkuHLkyD72Rl1vo2x44Wt5fRY1zJFybExMloLl
O7myGsb7T+E1NymwRANIfqRHmt1rFneNGUvsAih2QtGah8loX4gW7bZ4udacJL7C8XyyjWMch24V
mKMS9w21rOxYY2CORPgZ8aVr/8m8JEKpGEDLYoUj1YjHRFHU5x15Y30UsMb9wFPeg7suFBlnCI5t
dE9AV4oYFImbOmMIFVoWt4leXqsp/NivkuACdjPnWjHBK7tWOKyLrWt0p0mH8+wI2WbkWzDI3F5A
EZ2DZsnPim8fMtCBM4UXI4FwsIeyBecldS5VCaw5lRR0lhaap8ofTiKtyL39YEoRm+R6IqVCKtlU
rN6oRnXFoDQgCZhZPwqtfJ1lLe2uvFTY+A5KfHSs77kXStkvYSTRkkSOKyQJ2Mhly6OlnJpr0j1y
qhZV9GHTt65CEG2zJevpCbKIz6Sjn98fyN72PgXCTfCQymM8DnDrCZHcT/NNYptUEfEo6RewHj2f
6RsTOeHJaLJUxAaiMsFYSnN65y1GsGBRdAGB2ZIhNN4wejQQmu5rv0I9cm+8a6UiEeD1Py7q5KLg
ZMwNQfJ/WT4nbZKGIGXoUuplwMkl+1qV5h0xatrpo4RUYNSd2pdKAB7DguX27l+3JwtMfuIoyntE
0nALWjIMXMS6u0TGT5ieC+r5gsAE6Z0eMmLGqpvghGtNGRkNQclipqTMZkAvl6vCyzGkB1GOFAR/
/R7gFTMzmKCzKrr+lLiRIfYU6hEZvf+NYCUhzK2Zq/MasheLQu6BBqnLCBJhLG5e7YkOWgjyqj35
yt+4I7opDeqyLL7f/z4+1vUF/x8KFrFS6vIZgYjQmBnDp5aMQps96thstX2U0NUBMeuAVf3pNwNY
vkVVn5D+FxZwDMUuvQnvX8W/bjDiWqywZwhaGJfopkYrfJoMugseO1HlQtFXQB4u/lq26cfU+4iD
xo8ZbMVMAMV2gkbWxzG100t3mWssuzhW6XFXIZR8/WgdE2lZdIPKtrs3i3hcnI357Ytfef9lE52O
3J2OjlH3uGofpK7qp9kiZY0bdbIwJv77vt19fuMk49NH3KR39tLEhUlRo7GdAWjDiel1SRcHCkN/
y2x/wDhqJsF8X9os+pPby4aJh0Ewpocsv2lQ2g4oovtCw9V2rWWNFWLqx3uVwV0bBO3JUegVcYAe
acjUc6M75ukmz86Vsii6CZ2j8iXRBmMgNM0otj1FIH2W5P6wZyzTMfkx70j8uHJ3kD2CiwMmN3/v
0v4wY1HDFfwZa8N+hMsVk5JeU8qb1ae+m86mnwULWdTUGXMU85/V2IVJ0krLDnUADzyYc8ney0vr
iGHkQQHNbQ90HuWZiXejuFaxwJhI0Tim2fYS5eWQdmwbukhdYeCs4U1m93ldW5EIfOncPO5EDsZV
HhLEdCviOGkjzwCWKzeRBcMRdfampPglkFzarb8HWl1J+Af2neu1HHMx/Dy2wHZtkYfSi4Kv7vMm
2lJfPlUfbrBqAliALHQs/M0grO44J2nOoH3m6RdrpjKScZ8TapV8sATDxp1vGeI3f9zAgH+n5GrL
rGL2ncy8639Z2uTp8wWheYHM0GsYBLvMjpSCgPlPe39OsdYYEuuwn3sXBJyRxLnL4fIxVm6kd3Y4
XNxtZLLIA14yFZIVFOIiRuAG7JEWmKauUpIWEf3rysr+QXs+o1rWIqp2aizUj/307Uws5f0Pdh9u
b9ZFeF0Hoqa4EWLXIRzQLRfKymC10f/itP3JgfmkTv1ghbiM1Eo0Jhw5ymUulj3iCFL0wJ69R1B1
fqTsVdKo/CFKTmS8fKL81ZAnquaInYkUzmcCGHPFmSv5c5cpRiUQRbjc3xCIcPYQMivr+5E8jMfv
PICbVGKtx6lbZnHlya1fcbTM/yHEIQkv9vwyAjqX3luQ6JuRy1+H0lTR38mpZc9SN2EraGjKAuT7
LeihZ2vnn4BQMUqDmiFls3nq+7hQ5zp2atHjZpQ1M6R3r9vtP3lnW81vlWzf7Ovfs7zJjkAlVW9S
z/7USf8OVNb48TfmUhm6QDImr7RJrHOiJnZ8qKUAy2dvoJIMLa0ffb15TvvEUEA33kJEVtxszLI7
PMiOLsw5MiOBbs1SEwJ6RJYufQxNnsjMlS2KwF49SHKPdVXoW4Z0QqH/RZm5YtqZY85nQjLVzY++
z/R0KE7wYORMszNzHKf2P/RRqmrDN04n366Cha+PWdxbxzV2FvheS/BdPfJuvwdqlw8QebVmlXdz
H7DQB56wiRHd3EGwmQsgU0kKNP/YVHxEDJ8xxsGWbgQ3uVy8yEsk09Os/9qh6fHil65SZxDWHLa6
JT5iUshNTMzgBGACQAnxtGfwjT7p8K95ZDlJizj6dyzyupj5C2Sj3ZiRQdcz02+SBve/D3PsMk3A
R1FLYO+Jf/0Pm3r0glAigr/IajZTxM1rI+vvQUCWwJKmzGLEre5THN2w387QLKj4EtFBM31unCOx
fSGFCObNoTzcuLARNi1aeOemTV43CAARTeJx70r2r+al/JG4KyrTdnI5RBOn7a4zNEs5liPV8sB/
qITP48sBu4Fa8AodpdmT27fvbmnBJFN3MbS61k/uoSHwoM3DDpEjw3fa/vUwVjTVcG9xdtAajyd0
ZOdwvOLbgkIIEv7MV2U4+AdawadFBoc1JJgWGGaFh7kjLjrXAVDVejfEcuNLnaMBylOZRYGvVugJ
FUuuT4R2wGrZ75odKqhAbq/ri4lPhYfAmJhhIJR3MNZoXIdPvdSqff8sAPqL8D/+oxYjeaDnZmcX
/VrmpKhaoqPwuTMVfUh1dBcL05+8K0IVDgOq4ovu5v6M4c716x701zCz90dik+At4RLj5Dxb6XZd
tyNYkHHAsDzGI/HhZoTpMzqIZMdboXGq2K777BZdmxnVvP4+C5Uwr0N74JQZfU6CM8uw/oXQW5qS
/U0tODdEOgPiwFrfCJCHxLhWqcEXxnV7BwKSH5EF4n+85hT8L9o29epbpoPONycqWgRXNCgkMBPv
j4da8ib5OHMq2wglv4KTiOoRaRxTOEDkjNoqdVu2vkeCHDpsOJ95W5F5Sv0GIbUFHiaqOM+38kOX
RjTNp7Dcp1VsnDOao69inwyU0Po/rxBApfnwHBF3ISoqJ3+V0NMwjEJVypDa3hFGHupvOucNZgyG
U6N89sduFSzcq8wruM5dgIBEvf/mCHRtTCjapMKVEbWZS1yhisEc1T7nNRSHEZOLd3ZdqQL7myGp
HHNQJsHypoJHTKJqfS5RaX/gK0k821b2FpV/h2x0u36LFcsx5FbPuTUvUJL0VpN5jyy094YiFeky
2ctfeRW1zzCBOTvM4Ag3sEZtjcBzn571TBMHlYQPZkZOPJH73e2Ch3gL6+NQU9thXlkjq3qvqtGT
f43XeHN/D3zLnItGP+rzfJxdwcKWf9oDeunjEMefdovrr1j+uBSHtHWPLhSjvNJ2ZpNOVw/ADK7F
riwmKmtUn3TWE8ROJdBoNLWXQ+oYsewfDbPnd5BBzpcUQWskVWMVem4YCjXAoUvEgQxpdQUmjkwZ
67BCME4dJPMo/RX1Cv14kbeufWv0oWJ653UllyDS2CYFJKjBGhsAg9uaT3kQNBa9k2xE3SKJA7T3
DEWL9i8Th2P6qRbRSI39jJThJoFbDKsrgoFxRaT0o9bfiPsYtA1dfhEcy+zqKFrA7R0EDnJkTeEk
0D551EEiuGJzEHgCAMTDs5ABApZg3zdMyMvvyxM8nUSeYMJbDOd6Vh7nJMjSUHcwGoZ+ywnyqoxj
xM7KdhYGHT0h3u+1VhRa/kdQu6ZA/b+5Pm7+e+urRwlrmJ4uwb98kPqVtcIEigzfOEDphi/pHHTL
UifFd45sOFfrsQ4w/ut1jn2dY6458lmwWC7DfHdmmnb+M0q3dxvrHjk7tAlc0KMJ2zZf1ImsLn3O
JWPPaVO/k9OAHwkiqxKA0LPXbc7+WSemokg+UqECnJGIJSh51wqox87I0j0Cv4hIi/wi5O7DH6jR
hZLZmWYGqBp75hBZq03sndLQTyAUuqf7yNfv90t2Ej4Mj7JPpEat5v1d5sRiopLVU6etPCCLaoUV
RiM3Doiy+G5Z+pjwVP+BSTyxWV/MSS+kk/iL5sTodvlLGBN3wlE4jFvs/Hrv9n3k/KShox0lfg46
BxpKX1/t6OlX6rxJMdpRuT+f18oJwwX0rUCs4fX+viB8xVqIsK7z1SCkvOCuosnia5IrA3N43uq2
DMqFEE8gEmHTcRp1KXT1+f9ND452eH4WDGltCXT8RqQa1QVkeTEzxIG6u/SdERomgDM6HmTzbTUY
qFggpLiY+hUKjzcXJNvcAzFlCBs2cC64f1XE65fa0oObBjOK76Nt8yNKz/B2OCYYS72/8LohkeVI
3JT7h3HozHCAjvMRaHkbadJm8rjnCNcq4LKA1KPO17WIlwRO9ZfLsdxqO34Rc6TN1qp5ihiU9OSG
O6pz4N4CC+AJ1TBywjdpOeyw6fCu4+WHxEjMKR5yunz/II2QGbLT+Y4jkM8fP7lbSrAQdHj2ltyL
MAfRxhsNUIEYW0IUpdkzOjCgdZ9Jvi45VDlwVugW4mzzoq3LWmoAxM6EvVtlab1gNaFIBE3AcJDt
v2sP3YNJKtYL3lQOwhWRyc+QM2z8DecdhsjU/XpkLuNeFQjHSY+tcQupwC4C/xjRmJMxEuKK7Xaq
0e2tVi4sXY56BE3VQrMaN2xPPhZTmyXK8mBsn6QnxzEWf+axhaubtE03JPrvAJuQnUdQnpCJ4UVc
TuOTgIyBDnfGirWTa3hCJCrF2lEw+cW6da68tvFBhJiOPQmj1WyfIdqhZSYGEKqgN2li1YQixl5Y
d8TYvdPJxSlzEKuWW2e3jPhuF0pVhe9RWApPCMZK/SVN5w2oOzzbNHHTrba7bfQ/tm5ezRX/KaBv
teYyTZH5Xj3no7YIfi3MJzjPk+zsMMCztBf6bv2M2hNFtn5kVlZF1j4NPdOi5PzLfOMj40Tz7Gpy
goyp1gxPyLegnnT8Q0rjax369cbee5V+LJxAyp6IU2hVMVbDD83L0eARvXUKHkvMEZ8yXfD376/f
EgwcWdXRO3fc9w+2EEFVKBHJ/TJ7nYF5IEiOV9fbgTHzgQYGW9/fmNf98zK6JBFknD+WKSoSa/SS
d5JqX517HfVCg3Vxb1zl0jUKkfDBupcHRcUh7wi0jG9AWfIjLF+sbOrDFOx6DsSPrF+5wfdBCfEJ
p9jQgzOtlmzd7QBurVj1Tf9zJoqC+y2YgYr8FdXleeEP4d3Lm/w4CD5vju1mLkle970xhA6z0R2+
s/nSenCk3Ln/Dos4hdZtovaEEXKP9UiM7ce5FecyFVyQz96qjKgeHrFOZTlaLlcowAATeG77tAac
yyQYF/8wEUH7KFbeMUhnLEGHJ5LM5FGenQkWzPRRwO82xcWni7eLtBThGsZ4iJSg81unDsl5J4MA
BrPKoVFKgkrTAzD7MWks+rHKsXqcP/tCX3LqNEcKgDvUY6PKohLC0ZW9GLuWZIiZpvLUg0FFGSXw
wOGuk9nrqnBnMAvFviYU4mEvzZxaRuL472ePhpYJ309Bp/PnNSOVpZwbh0xUy1O4+aTFP4WHqYBr
68trPwSl+LrYQ44rHRgrne1kadwrT5elEW0O19gUcmnPbqaF/FwmtWW9O47Vx4LXyFT7bemM8Lif
Nzc8Y8qlZNke4WlxHxuRDZDjJI1IM75OMRqHy6gQSLvmp/b5JZX+C4iM7eRCWtnSEtGuYMFFQKnW
nQfOMGjr91eEJt8r6k7z7LLV6UGZ3E+/0QFPDvfvwuVXxObdDp5yS+QAKAmFA2gaBaCbx4wiPTIV
sSHeDzgS3hi402cfiuHwHlrZ4oFGxL6iFkwW4dUNtdELZNtsLoBBhJGvKmHqk+YihURgF236ie7o
OA+6PY3eVAcq8QeeFz/lisQl7QKjVKfUcZ5WGZ5SxERmFgKUFSc7oyUsZrQSCAYK09XJy9yfMkd/
Vv/xH76XKO5L9axjxcjObtJQeyKd5M/AV4n4NygeMiLRMYUyFyqXVPkZSeTZsZmVHhdCAb4x0Rdg
SbiM+mLX3QU8GTJU04fBqY0DhNh9vziQFsU5RB6OQZD764QWaPi+7ceSnr7LNiOHd90ozeAxUjtH
MFPXVkgX0VCuJsAiRX1pWJMJMhg7gWLsnGrd/L+E4BYpWW7iX/mZJUn8lTiEvnbreShyMpEvLmpd
qI+aApiteTJB1VWB5HbddYtafKA9AdW0zk2lz8XpN8RxrxM6xCtS05gzefeteclhaBRov6tSt6t6
kpDw3IVVl6lAENrnNthErYmvKKxqfB4ShVtpVM7Q4CYg/YKHrO0wFcbuy668j9VQ6YBhywFpynbK
9XYvJp2yc18SZnsmtNfhSHQuLxpIDVI8T0GEZQYZ1pF6q4+dtWtwxTDv83gWeIcOYU9Cwef8VisU
lR5/kfsNog3zx13UFNRgJv2d9huw5YxVjZaV+VPPgfcYyspDctDMqGKWb7ursqhAGBnEEjgfAqoH
QfBJt+e6w41SKjv91lGT7WcahpqcMy3hYv0OYkfBjqROFWsksUSgrdfJwVhBkui0emyoi366iBOD
nGuRsASQp2S6oFqBn9GpBiv51UaoWb5hdFUSSs7Fxj9fkYYM44y121SMpy7SvZ0t6zeor1gJENJI
RdTxIQHB/riuKzevaV6JdjzWSQb1YzDC4M1iwkuRmM+WzYLtDXglPKIqn40xF5iKLB96Xv1ydqts
zEE5DgYFmWPYVzMcA7hDogVRnOjKnrNe9ZF0tfqsmSE/0nUNQCiwm+5Sh4ZrrwSmWYxq5KB26uhq
Vk0DQPM3kpyES0rT4BWPrHsI1w+EFzdvODKafWaWdF+kcybkChENXxyCNy4TkcHuuamzQ/ZYLqLa
gRsBICWYZRdepbos0TmwoNQ4FdYRLCFCI2HFkGVqNEXJ0AwKN3tY3MAiTM3XnUDulSHGtHRRR3Rw
tCcgAQsOaSRlBBHkTTOTJAcKcehoXZrTlpfvEEEw4PxiYFGgwM2wZ0cElYQA12xHUMT4AiaiL40k
TsLXdDtPN36zsxgKCXDfihE3RfgaKGDeMgrp8eD02iVZizbkjkFY2vcL1AN/KXDqhIkvR6UDr2to
e7Y/TnjsH5Af2+1prB6/wDTsmt87cKmLgZDfnDOloM44ZyBbfsJLNcBKjODYQU6A2HDFykF/FaV+
h8C3uBiNbQlu3+4OHhEhuZa5UZ3C1uWmR0LuXqjvUQcFa9h07MFVlG6KAoomB2hAWU2sbi8xx4k4
jgYiza5DVR5LrjgqkbNKsHYOczQ4QemrrFvFcc67UZqAmIc4dqvVX2R1nmielPfiB/VkBdvaCf8k
aOpi5q4BeJIftYr/oemAaPGOhNZCD29B/NXNNS31dfHt/nt4E2rCWR6+MJV+RQQ2GgsdYpv+qgXC
kcCDpk+NXd5nVsmDkJRJ58APg9COlNg3+ih25PhmpTLtSc57oyqxhurjzWzrMVmO4++2U1pE32Gp
isIf9jM5OOl+kcflkQi2gq5Mi/e56aZNDeWroxig6FMP05E6thkR8HRL6YPMdMET1nCQRzFuZUiE
yLLNgD1alF/zdYLe47zyJWXLivfOeo9XogRy3FwaO66e4zfyawus+ywGdOFiELb0ND5pE6B/q5b8
7iPKbsfTJqMkf97F1+8T0joGyVbAfdiL7rmwHItF2lnvyUWt7ycWv14ATOzuCBP17GvYbVMAsi6X
6SeGjLK74Xnftc3pCSxdGTF5/1QKFUL521ievL2MJnDQ1YYiae3fULG5RicVDeDz0EY4jG2OfkYI
1zcERpJhL0y6hfD4Na+/ODaPjWKCoh81/Hjd6MRlZsNo+MOL7A0HUGa6GCG2sN3aVVQGttKvLr5H
ve4z+MFy1SfPxJ+9yQHw6qeGWQOacACrah8/VjYUvzXxVto7jwTaBkGsZ7MbX8CXwl7XTGx76M+u
5GuLC/ey2EXLG7qF8Ipq/Yj4ANzSp+50mu1MF8qoTGundXWWY3h0xn4Ul0Mg39ufCX3K1s0hUAcu
HaSJqd7U06Vi0M4FaEdd/QEa5IhE+GS+tyw+AZJAKOvMcnRFhYPOeIi84BgXpj9KsyovK32OHJKA
B+9CJCjHYCponGodz74dpc3/QBn8a31nlXjZO8k+9yI81CTdHQrxzF94Q2gcFcf/ep+Jewaf3puP
TOXHl5ueW3lVE8T1u04qYXJaBsLAvJwQicJvk2PktfudbEX9N+0+H/1nkos3odEGd10SFBMgBFni
7ccttQo+FynFdkgyqA4Bwku/fNUDkIoc3TiUeFrlnH18gAbHn84OdBZeVimHkThUt/xYochLZPAt
njShJBAo2ufbkrDOLXiiLn8YRUigz6RAnbbaqfU9fUPGm+3rIJ/7TJXSfCJK+e9BGRMzHXSdwUd1
dedwS1V647Lhd/tCGn/Typwu5x2jjGSMf3kklv2yI2SzcobiVcNmzzpF6dgt2mVBBlg1yq9Vi5uT
sXEhumhHHhnIbaS2TVy/B5jsHjtQzUwPBBvMhtcoHCFs/kct3xBq9R9eZFsXHJNZTz8G8tlwJAq2
5+1Z90e2mFhF8RlPL2VgnEMVVwnFhrV/TlbzDxxEp7p9CXrqBcghJbUEgszehmhp1WHbZb30Nxks
TtRkMxKRI5d6VN5zx/FUszoBsjVL5MgeeUcdsuP6X5XihD8WJlgahX0+j2cIOTHZCHNbCN4SHaVk
/V4ultdY0woit5pF5w5llIxCpvNLdeusV+Bzo8HaPAGRT8hUyn0mC3PVcc5N+gKvMjb8Phxvdtw7
KOIStTANuFbb/EA/3hy+Tgz0h8ODVn4Avww9tB7YgH043LubFmR83D+w3f8QVRqZz1Z0/4lJjU8c
xNSRwqGBs0+eV6nd7pYAsGmJWd3cal/mTQhzs5fp1v9zcaprzFxcwxeUJuXSglMI+9jAfysJUbOX
8kOcAyxsM5xYq9OrBN1KRnblMoGW35iaRsHkSl14PKxvhQuOBobFZaOts6iJ0bZkk+mWcdLt12e2
MnJHkK8jSe0BkMPTj5e4gw3uecD5fWSeixmFqg+swyIoccQLb6LusUDjXwMped5fN/tUWG9nUljT
5wz9xom1oAMDhMcghT0SGJrTGme5APl4CS31eobPe+MrVAUVzrgZggoju0kEi2PIkgj3//JskqSU
WmlFogsD6swfvn5QqmpOU/OfNei54wGuguHP2ZsOt3vL3vbmM+jGNM5ubG6cMzylhdmEdaEmEIqd
muwCATI6ZY5ZSZsAd/jHnJqdhc14KjiUwLvSKnQEdtQEL0HTyQQ0/A9jJwAI/7IcWGS7FSFyXpjG
T7oRt7+ip6fYRW+0iBis0WvGAF2/XwCFbRpKOc1K1JfqXhLz7YNrjojnGjI+iSLtdMGhMR4ukyc1
7dnm71kvh/GGJd6FTWwCrS03DAdjMw1LUMW/IHDsqm/YlYCj1Q9EgRVKisc9gmcbFhmk4qUXPnBr
xtGkhi9Y8xlwRsNLmdoHfQjBjK7KEyFBpdzzR8DuOQUUpdYZjr3NbQWrTtT3KzWcdZ2O7mnuU5fj
1G/bbdOAgQEqpTYIBVkyjaWZGcKu3hSSHlWqgBw7u6MCDns+tiPD230Qts3ZxAmsSC3xbpf+0LO/
UilPpjWWZxdooz0fAM2fdSYBYnKLJG4AJedpFPmsQJH5yFkwaCbhxHJAzgdZbjAlUo4OSXg0Sfer
txBOq69sUrEkZEmZyCQmw6/GAJTASPm8ih6blUVwPYD2zNptpl+86Xg0Y6qpLsUTdNeVwRseYVhO
P3+cjzu+qjlA+bCB8pTPRIPS7PpfmjZRXWtkCCErPr4KVWllGWdZJKiaTkc+HLJx9CHstxUJNyVS
Kf+fvNPMpb+3LCY/t1Jee+lq+SRkkhKSSii9GY/qbB6x4iW7FIA5bQa9l8e+jbBzNhPYXv8uvQmj
4kvRVeqquj7YsddOyH6lhiPP6hI8EG89i5usJhh8jSh9mJRBefEX3XwKmKiDbnKmpDIxCpyXp9VX
XnNmMdoPRXKmnoEFmZvxkEls/ZhfYuWhwZ5wLOSVSXdURnbb57aMLylFTgxpCft6f6/BbhbzTB/i
pLTkEyxeJQSIk+DDLpR4s/Jk8unF5oT8+ZJAeX3MqCv+h8yosG0beLnLOEptP3Fpp1luXf+bH2Vn
nDjOLXjZMUTf6HYafL0JeyXxP4oEfSIIXb3sPtx4EeZgzlOxhdxNepFt6TOHEDabh3tFesBRtc94
RYaBx3coNuXRhWEPRi7xi76CguFJjK4XaClptgvE0rczz44KNgmZfF8XSuvbR4piMeVMqYBh4dew
NRNm2gLTGjP6spWKjAtrCC7bQizx4sqm2aRiniEuhSZHEHf3/q/sZRW/0NC3WzQDaa+pMMwqjrT4
WM6lnJUCE8BUlmocxai+++UJGC9EdPzW3UHdrjKm0Rh8fxCse3BVl0WOqTHdWx2p/aeIz9hyY8hd
lmSvb7t3twOUo/bavB5y1Rcg6nRNrPOP5aFZvA/qqJGdtuIDDr/G0aoxVWtaDxDIENhs3UO2Lgfp
a3BBipX1jM0oolQsWg+hIu2jX0cXue1XZVQul3Jy8N0WKPvQgkZVgIx3dMG4UBTS2jOqpMuZt//4
r/dbsGIRS/JZJ9Y+XjXpqJwnV8dDaZ9gHHbF9pEY4riZZdZfZFcPJxu9faqNr7Qb4jOjeZAjK04x
HcVFStMUTOZotUkf723Z3soyCPdUi203zTfJk2mAiEP0Uf0ezGTAne0DjLVpAFyuEzyR3xu2nxag
nDtwJL+SY5CtHguXWZMan2bGEB55kSE8eeUE/0auB+hZRrdLHLkJvvqvsUTk4n0P3vlj3hSw8gaR
z1kmiKvUUGNCZIcpVnFFyRfkgPYCU7uxh0WAg6jHgY1SqGHJzEdvAKpmtHLkP8zvfiLccThlWSTz
2rRlDlUYWPTdcfg6E8NZUnH1OvoOp0bbuPLbGB4xggmtfpvltiHChTNdFqa8WT4AwOqXzFvNHAPm
kWPrdZ92wmtT5xVK2YomfAcfwllFMvznYVJJ7ihdD4ZpvTJJkohuwjLGTStgKRmOlwDnflmF4eSU
ScUMaSIXA+Iers1E/3gXjS49P/MGkEQCRjjAEzOfRlA2QmGemQyUfnxXTw8ggviXvkfxDVdyvxRB
nY7ZKOEsF9JEpmRHx6BDarW960AEaVzJq6hNdxlF+1o2L408MZAPUD+1S0LS7KO2mdh2txvD5wil
HWIiouS6G72dHBCXyU5LuOTlKU32vk21Qkr31azn391oRMsa9SFBkFN0jBdPiZBAYmx+RnDKizAF
S5CXF/j23SepaCD3G2yes5Zibw4SZPwlCVd951Xe0XmYzDacJdhMYTxYf4nBzNzvKAS9fGVudG2F
9Qfeeira65lU7UuSeq67NVFSh5/VvAlv3P7mglOrbfnmWqJlhUlLbhC/VB/tpvOcmPYbIZ83URjv
YEnPEXs0DVmwjYQM9kVWVcTRZtl65dPflSl3IjThHlT8pq3roCHYmgUjlXT3KjCzwZ+6Holrv5Tf
/2BxkOTYmzPbeUr/zl8KGoSo2TVctNZl9Zi3beMcoIk7G/02Kx2VwtHQKcz9J3tXzsWFf9zUCwTf
wFCAi5KS03rJATxP+MDIGRw9BD4N5MMskaPFuxUm/x9STZw0nfgxWq0YuvW67hXM6wIWrgdlnBUJ
/GBLuRBNGhjYXcE83BQwZrQbxGeDnDX4zsHqOZZsB4DrOlfqiIWaHA5lZ/PkmPMIUpg5Y3E6XuCe
SYQ3mj/QevYCoSSVw4SZZsunxnDG/0yh23m5FMKUy5itoGri6/7667Zm1dxbMyfTcjf0TE4kfyJp
iylJT7XKc/T8rvshejuZJ02G8M71wKr912s2C5bUEP5xH+oPKiIB9QMifRrehK9v1g6aaAWW/96p
k+1qChWkCWQSwhjpZDO2n5NltXupsCL491UYWPwUuQ5uOlt9jA8L9dASTohi8m0ntFhQzGRzBI+q
/f8poyLC3ZOHuTWWthjJCfe90SWoZWO7JawDZV7hi4I+FkTrSsheVayvHLCqz64z8B1YgZQihnAD
zKzx6Jo/+KWn0KzWAVZKk0quNNLakxksUZljH+hO5M9wLG46JaLYo4ZZy9t/wi0/AkjeiNEYRQ2y
PoyX7LJiNyDxI2CuoMbrHdKtCzTcEk7U6xVESeB7jEHiavhmmSDqYod4z6f1rNQUlIxrcbjXD5jJ
AVqXpYQYSIgxgv5BAJP2srNQqMew+T6cec37lfKYbbQuAGk/aXgdDG337ORioyzWEQU2UL/UVrLL
eZCZGRp5/tKAneN2V4XP3Ub8YlwEa7Uu0ej6FVPgQAKrvGARAsdKJUo+VVQoNh/chuq5NoLQXiHK
PsCH719AMnNwQzn2t1y1hoD4uR+MYxIYPmqBqovTtrWeMifvV7DE0hpEhfLkXvhR+eeN2wrWvJdu
eex3Fgv+ndrDFGkDS+jj7jESiIqywL4XvXahi48JLyg5H9UlmV+NkxoDRFOlrg/OkJ48iIqAnIKN
YZuXJjahX7sgITcSD4A5fxSaocHxua0yd7YTkEsXbPBDKi98YM1SlUv4VRPk8v/E9FZQW4XIRkh9
iY0pz2brMPaB1Ps+2aVvf4YPo5UEqyqON1C7t0dSXnhMZdOe5pbEG9mhJynmqAIvX5YZ8HwJPTKv
+7QhpfaeObv5ZN7jallHNpb/SVSJrMeCMiTcIHqiO98gFi5f6z9/4hUWKC0XxLuHUHDC93tP2KlD
BLiNQ0mX2pjdjfTk5v/Lvpqx30HGX867VLNVs5A219qlSsIIyn/RH8ryAAMcnA86akCFQeE6Vvu9
XAL+WSqLrqNSLFvBqUTuC2BiDd1oZgFcYyR0lqMEkCTFV3h1KvtHwcBSWLXO/5IotVCkJoEhDvkT
sAX0cN12n8k14wn8Tv+nP7yKWofSP4ydn18TUx0necB2puB6Wa+kqEGEjNytuzdWKhsyihPRCwEK
wmU96KuNcOpHjfuRN06sXMGw/3T3h5/ZUClurjrGuRNMRjk5dK7ANHEz/+BrNpdq1liiJ2qHm0qt
Y3tnUEuy3m4o2lo+BsMNqltXeH0ltwVPhdKQjbXmWFqu5hwRTL3Ymf7M2p2/ZMIcc/VfNw7Skk7o
12/cYvFhQ0oIl91JNpsYr9KRfJck6xE38kYEiQ+T9AawVDxNrkDym1Kz714nKffjF4U0PgF2duLd
nD8j2fM4xmY5kwdGuhvGfKz7LLQ2nDtqR1UsrlmoPlI6/a32duEGvww5+U64JBhoEH+QmqnMEJKX
hf9IeP/muCKPgvV1fNRtMqQg84F8ZgDbKaXeP4dtViXjyxWjFX2rYh1nMcY/q/GS4HD4CYOvNVHu
sqUizRmpVG/NQ1yxyJ0RJGfhYV7pPXIvtq82QdBvoCK6FKi+rWZ6RbGvf8Caz3HT+cHhgs0RZFoL
ed4qB7mKa6Ze3pzxxJ1x5T2zGHYz6fYmK83cF4KuQeODvvcqv6ckCjpmH8TV3OuH6W8XzMrBUtzL
q76RSffhniPx5aqWEBs+dlqtf0WcuouCxyf0jDLeG7xzJQ7Fc4ID/PY0tfL5/C0KJKdxpo+dUfMy
Df98K2j+yCDbpbDGMiS47AUb7q+G1Mqr+2cDRhcXCHIeBmwy+UdcygkEPK2nzmb3VMesk+cLOo+Q
JMEDppXuXykccbetA6dtZ3y+uPteBxfXizm4hm/yU4n0a8ZsKc95H12yUz+d0Uzm6IN45kmhEFIU
hxdFv+Ony2eNfpgxafzLCnngggxQ520Y5kePEt+yQNtO1WQWsefyZt7MfH1W9cdOmoX0HfBcvvsF
9q3yc70ZBriRbixz/QSCb7OwZxopH719h2hvUTh0+MQxz+pNiIBfreyGIokjF1jX8vk0ZVR04cbC
K7ummIvAnsQZZs9g1faRyUw4LDLzSa+evItPhh1D3isJEK1X0VjCDFLT7EZFAcsG+ivyQmE9+s25
tkQsHk3BbQoHfwYFLfXDJg91ej8drlEx+uipZp2Yde6RSC5ec45aWICyeplFGesBvWsOYJYUGAoC
Rd/628D0q6rhcPVUrG1f8++Yz3F3740YSxTS9bXsg6nfshdq1YY/LnnP6siV7cAYCdpJbzM+WnUv
cOGS2nPvyq30j+6TF15bvr3OCg9PzJBnwtavTbDrybrnKQcyU2dZFWdPEFOkNPVreDRrtiL7Qn0k
TBj3GPvyhuSu+8aAttCMxIsvHxH3ZIQpzhDz8RirxguszIZYdejn3fuaYLyi9MO6DzebsQ/NsSpY
3UmgUPrB8rJyCgbuGvWQoSfGw5N1mAqPklFki+bhhmoF5Xfc58wIt/dv0M0lACcMg0zYDrWEfAh8
lPUmDmkjRTXA006lM5TNSvfYe4uWzJWg04FyDhKiR2LGC7pTTHcd2lsNTk4VorUnZxMzzfJfgKKM
0uWzIbKcnm2UGCpNsmYhkk3u6L9Se5H0L2xiAn5+WfRNEkZRbmE4pAGohuKJXMhUciX9TGlWm3Fa
NddkFZ7b7tk1/fDbCd6SkT881Tm9awRJyySMr9E70RisqIy+/Xxiy35X5kV2ZfvT46zjLCvLljH1
Ab1aYeATa8g0HUPPBLZwIBSUjz9rcyb3dbwOf06hhPYNS0sNdK/jixFNaE0uf3DTqHMOkuFUZK9b
1pF4SDNLw2SpXvFFSsA5aR9kLfkM91lOZAEC2MLA6pxkfo4p6XRf6+hMKDzligBlCFv4RYD5poHl
v3dka/DUf34xnhruClRJ4DQGFAo99vIA5aNtR29gAOcrLh3xYtvP83PQOd8qv1M9PCaVQF+Ybwph
bEQ99jGfeNheNtewFPLXKbRen2WQm/vWX9nbk8tGjvBZwu0drXH84v5EPOiqAU+LFIWHEnE7bZVI
q1nooAsv9ZjdfYUFB/1AHUTRKUKifSlYB4o99OzN8GLqOTGVXA4oN8mAv5fr44hwR4mQY/4ACnfz
tUyWfGcc63usWMAnJn9zZJC6rKeApfWhbcQ2FQCrOgmTDrkbm2sU3OXh5nKJa7dUNEahyDLi4TYl
c6b17GZDaup0h4O02ipMdohxjHi80godMfE3bAace8BP2C2uLqUekpmUACnZJoFHZv8JJwv5wnFt
G7IGFQp26lirAcuz4YyH/S6EF4C0jafD2etVwlUYd7G9WYd7/OujLH/MqWhS7F/GLMgydYnGLGNw
5ms2VZ3KjdFfY/DRGUGOscm9Lkra81G3O8/Kt2cJe45+xENipdnKE3nQSK04YoD3jUER0OvPtup5
WNzL9LAVXYlrXKJ7kfO4/refESeZolgUJ3rJ0K/gGN9Ilgk711MMzwtkUMWb/55BvlkPXTOM0BVY
R8W3Geo3/GQe6p9dTP9ZyD0KZBJPW7o9PE6yvpa5XuxFPaR7z92eDfWSU9S4rW4KEIolwtpVRM8E
Okix2YFa2WV1wuivmo4L7kPVykVXksm34WOlxm06SQHUlNGieWAFFHCAnK0LUHrp+HgKswuGxaig
G2H40u21V8oNpNnKhPL06Yx9mv7lzJ49nt+HwW72E6Iy2eVB3eMimR25WiO8u9KCoDnrxhtKR96X
aY6Ox+LnrdTmT9N4iu36jZl63oAXV4p7hFOX9T+HVqrkEUS/yXx6xA9JeC0GHJVLuXGfp0CV8ueh
gOF7VxfjStN0blobLaB5vWMFZuwdqXQtUyCwlRwljs7+6tQUjhV4runGJZaYYKrxjt6Ke7OkTP2S
F5JT7iwtkTTshyY5szOYrbAu5DOVnS1ALBhPgovKy0qB9HtUdJq8+CdH5YDglMQqowU8tFz5gacq
pedgCFcZEMhrfYYfcYicGG0BSm9awtdUY8xcHoaS7A+KXEa1HMSqH+usXq4cuvna0DgqlKjmN1ij
Ye1eLTcHsVpXe10ibFSEtaauGHF/QudnFpgJeJ8wtOn5F95mR/qUUJV8o++rEb/sQUJ7ZzQ9NiF0
Fge8cGHmzp3fadPjtq80WAjeJTgxepHo0+iEBm263o9KY5myAmmuolPcy2BkzEKmxdf6Qk+xJ765
ylCWHln2ilSPkqPgyqs98ywwK/aX+8TeG9lwptKOXnGnPmlpt02+5hiVy72NUBRD9M26OjwrQyv9
QbnIi2TTic/vcnYg2A7nbfBCAgBBw9FBoXnRxTSTFkBAZWHh2C0pMw2pGVMuwVN8Na5tscYsgBF/
6u0sYgR4mpvNkEuQSMey1T+biBi270XViqPiKoYwoJwdIVrGB1suvB9APkkFC6p00tvVNBCvqYDr
VfjkraLUTwmUe+pVrUDbiSo5sTX5rWmx8Cc2xPkbFHWwy79i+MzOmQaLf3UfMI2s2ommXkov3bOI
H/7ILfR66ImvAvBOPaYA9gXgvpWpqoqs//8rNIKmCpKKmLXMdZTHKtbM3NNvwkQtN03TPt6lWKlb
GIFwwRqJTZLwOHJEQL3WUmsUTibxX5YHsWBOLR06in4NrW5NvddjjmcLcWBbkJxb+8Gddp0R0vWU
deW1ppNE1EwCHZcwGZcnvZBuThRjqHzH71uwu7c6jpxc/WnGdDpUhSQVBxUJzkSv3cHsFRkuQNHB
OTTdFy8voeYDC5rCQGE8rLi4oOVtot9yy4KYBs1Amw3txENNsgqCcxCp62yasvUrxWkXGsu3onAh
N+8MQoXjJqVrGkxM4axDZwA8vB6SaHNQ8QFrwBddYO36bYX7CkDFk2OH8a0mJOcMELjnm0hqu+k4
w/2VjEIzrx7GYoMJUYDu0MC9jf2kmxzLyjocTz6kvud8HSskyV93IjExg7qSiBMSee/6RsZP1lkk
nl43W5R2XrYdAytbyJirmsdQrLAEDdB/+BxeKmw5SRmXuYHJPf7tPEtokwkGXOPHVYkjERqadPD8
4tB0h0565YJ1PxVZPbnKhoc25qabO1G0eolK5V7wl5wM6g+eNjm1QOE1r/Jx/q96TI7hHpc6wTnT
hZK/u2jd57BdcBeWhudmgoBoEM6bxOX+B8hctpmHqsz73XJEE6aPxdWt6/TiNYEsFJGpHfY98slB
dfEG8vPjMLA6MpdDGsWZ26mB2gYnBhMTUsUs1wm+11+yhHCCXIWBiU11NbpPRTmeZn5DF1DwLBG/
Yvj/Xe7s4an9hpEPAeUguqJnP40cQSkQyY0HXOCBcA3OKbwAhYPrxOTCq90S6pjBOSL1055IvkVv
twCPraiOo9qjf+rO01Kjm0b6H2qd26YiS8bwpmqg9sWK3XVGQYPZ21l21qyPBkeUC5aN20piuvQb
GguxHwRGJ59yLS1tFvhd7PZ4p9MkkpzyHeKumm4qZLMKSE46XuOyTGTEVH5R6+DoBWTe+6bOzktX
iPdX5u+7ltmpp4Xaj86wSmgXdQmke4zl9DcVT2zeEYmXM488+hYIY6207fn4TMhZ/cyMCNhI5Qv4
jFDUSWiIviHhsOuvVonIXb0k9SSkF1+eCt9PxsZNq9OgTDg8K4nIj6O3j3V7aG8wJqqjXZAh8pBN
AvqGW+1lGgu+wFy/m1p8+7IfTppUwaGAMO28TE8rWSK+d5ysVZxI81rtlRq0cuqxz25fgKqxFIkL
RjzYBimyegfSIxy6U17e9l4RIMBqiL7j81rQrBXIg8r9mDbW/70XrvDU/4+9Q8XE/8kUeepKTsM/
3qGyRcDhxxfYXcel0/qBaUX0z7KVLEO3qMOl9JNKEtZUjvXqkLG5k3ni3Qf/OIZDoy9isICgaBwd
zV97GMXBRinQBXWp9lJmCOzeUr1Idgcp485AJTXAEezS9Mf7TokAgosMTNN0PBU5QHNuiNmFPHD6
ulctoD7d8PnnRMDjI6z0UYeeGHP/BjV2GnyCq8qFyeZzohpbq/k21HhEJ9rkzRlUSo8IKk0upZTF
dAbZhoLfyWO65MKlKcvhZ0+GLZKSwHFhRcOhJ4DblAGlpLfXJlXmESmSn6D+CioJ0nvImvkVk1U+
6mzqY4Cgd/D3AnRrl4kUXstqU/c7n4RWUs2rPTG0MXY1AgNYhz7JJGqclLn5aRm7swNAVasd96Pb
A9a3qctGiOk6JMKUm/9BDbplO4cdxJZ7ZF7gAcWasjRJZgNVxb4AGIQfHhHXMbtWE2wexmKcj1mS
Q/CqWoGwzjIus2FLyqPu8quMgfmjjjJGbURUbJdbXo/shVhWRGlRU9iPfl6jLJ5nHiGth+xSnOdt
iuVJQXdXelgIBVKgNb+k/A+oEAWYVoxIsNmFW+xYGZG6yap+hYmi3ue7GDgD7b/wpUZuJq4IXB15
bVFFapXeN7h5rxkzSjhET3X0HIdVl32ShhlPKtpDg+eZjtwkrJzHWlbv3ayv0mOEYWFWM2e4rUY8
dLnWDc6sP6kOP6QrXC8nW94TVpwha5HJBM7r9aw1i+NoHIXjfWVRTx/R6SbmfHNqgq0MMNNyn7lS
T3l4Sc27Mbn+wRJuEuuMm8qvdWsIrdLhkR4I+ITPTN0JHMmkalcGc2drHGi+L9Kb2RJFpZA2bYJE
ndpSjPq08wDSGNBv8ZJm2Os2Q2mU+lE3gTyl++QYPZWWAPWf6KNfRzD5rJmOpDxl/ZXpqhjPVUZ3
mQAkji7Kh7JjkvXrEjXoOlLs0RwLgwlUoiJmui96g4XrYJwkjZlhZbanXfNBIY//w9anv3jph9gg
5mrLHcfmeWw+xh6Wwh6/8NyX+Wzr6BZhsphHvTQFE1JoYzZzg90NkgythjrH69PyQYaeUHPyXmJt
mjA0G2X1tzHQ3h6YFHsTiXTvH0jUsHjjUJW0vCJwHPN2ZGGkIp68B1jLlGrwpFR2cdQoHNv+LRX7
ZhiLwRQQFoaoKeShywMDf6goG+8KId5CzjxlUJr3McfjhBkg6rhPYzVlBAAYFjhdiselr1FoZhxD
6KCBm983J7Zksb6iQ5Wid0GW7RSW0n7x2IYS2V2jYfQAORD8QgaBm95FoL4qU6FA5SvRApSNZW2I
OLEkpdIk6c8BM76k7DtctPJp0jnt5UwDnBuuqn8raUNPb6yBzk/Bzvc02MyePibUDmh34cr2+Kcf
ywGSHLqT0VecrYW0vb5XUqbL84uyCNpAMDV5XGxQ1rjBBAynJcl+kTSKP57kzG96pX0osvNvkhva
kLUx3PT5SraDdCykoBlh1MiVqMtcxz52Bg+XFaa10QO0wEbBYzQTxAODyv2RJoasvZsFnN3FFYGr
e5VrWq5+IYzcXF/tUUEqy+RxEP8mmkylbIzQcRWwmchF8FkyGs1CeUjN6N2G+l65S7xx1BeGQgrP
n33bq9+qnJTrjkE4dPniI01BWPZ7FU/bo5q7lrl+90UbhNSsYxww0jGvO7S7jCLiwc+iUyGUa00Y
kwpDhCE9/RXHri3kk5ceQY9WxiLhlDZZeiR3hpiWYk+59MqFaLzzqunIFDLmrIYJkomu4UKMECwW
NJHyn2R8Zr9sUZzBlpqAvh+Q5ZtvT0YJMm0bwc32DsK3n6dViYowS46VPojFOot4szOhwH4aMEGl
3RXsH7bPkXhfD6xuNAafz3+AxJDuLuclJPdgMGjaL6ifWCPKXejgtQW0d797g3W1ij3WixH1a382
ggyXizBZQuJImp1/Hd2BHVx/cG/9UxYpeQWjFKj0ha2W1MksbxUOFqnkyAMUSkVnUYmwsjo/Y3fc
CKRkAI/9oMIk7mte0aHqiKBIBX/RNrMRgI2e3NdPExgI/UZO1zhKLpp1ds6IaerdYmzpZ8VbhvHH
HcwS/jR0S1sZIrZ9ab95gFnHzhCzNk9yKW4V33+ONZrUFqfitmF4SUZU2LmozLQ1Pfh1T7p0howR
QPHGkYVRplaZ8b0FXlrYrXF/eazGIOvjzRCRjaPbUYVaX86WArf6i7DdHXbCTOGGeFyr6O9bMX7j
inzz6O0npWgQ6A7jNmMaVX8kmI/R/j1nZjtZ7lGnPXaz84Yrl0P+ARpH3plzniu9n3o7pwor5y3a
viTk2lu9wD5rytF9CYWS0x8vsqYIUOiGLt5flyXHScDxHdXoPtNOVD4eNL2q2T7szDsrdhHkQzHK
3rq2NCXQoELwVIYMYrJeiwsERRuUIna8oVmVUr7jKZ4Nzu1vyP6fKVzaKHx/WMILzNfViC2094ul
FE6orqHPxTfAksVXhPcsAeHlY9K/Iz+wGHid6VR4Bt9Unzt/TrdmaHFVGnNIMwSCAJjWzQegw+3T
9xKny/r/Z7Fu3fL14vRJmm81BN0c/fsasBGhacm0bP3xBQGvZ3Y18hpYUYRf421NgM12c/9XRJh7
vArjSf/RJMwtfnXHUXliiytilDWy+n8b5wcVKVSlE1UxoZxjhqWWV7FK38WbQnW0UT3ipj648jXy
Br+eHVhlyRrS8tV4slFkxfM383asdnV3AVk4DstOZUGmUqpXZTIiDxrx1no+SQXrhwms7RwoLAUI
XFSnqmrccm3jbnlLGHbpY0y8k2pJrunBIq3b7RpCTspJCKdQO6OsaPQblAOrebSqJObc+xbGU8Lm
NDeh5mEEVy3/traOtE1OK07e/4qZdtWnZtsC5GWkAFboFGtlYrRT09mv5fXnyQDmwuWweKwbJZqA
hpDMYnZJrMDSh4cTXrUWLoSpSE92d0ZkGzMXvpjwZfkkpkS7ES3swXodsR3Wb6iJN7r5qFMplT3c
W+68iB/jv6b3I9Tjr1O739pGFQMGeYkAbeaNMqCX60BgScc4bwfgTjIcBtMXmY2uLrp1cvxe4w10
L8+sqrM9HVpiWR7Bz1jtcXgeaw7YpzMr553ZJDl7fFtHrlly8NNncaWB/hF65zk4QBqJg4f4Tt0g
IJhTVpXbQJoIFKqks9ptOFjMQt6NWnYwCkSFG5rmFCRDiFle82e2MPtguqhjYncjFqWPaPcVHWJB
YjoCfIivA8lLRL+rc5yRptVnHlLe2/r5YIDe/f6+89QJ4M7QwqDQuKvh6VfvlCIY9UZu4FwSaRWm
osZF0MEt/ziJyWefB7XXOhCXFfbpEgnUKbX6YLwld99EP/FlDDSM8LRQ7ZlB9iGAem+AizbNB6Fx
Vy4tmPeKsl8vRdyBbHBgcPltVWcVG8ykrjk9V79/FawAe3nGq42Dm4znHm2BEloWWDuf4yNzbYR9
qmXxXxDRJebW7noKsSsbzMhEzdSk2wsWJdIi7B9gStPoeg+1EPlpxIqrOudKFFuMnaOybGa3Xw04
uOYtCkxfrx00ggwNc0JgpGdWLMc+pTUo/xtvtHtRtg7DsB7aXa/dZPzpjVzc79fOdSz/+1u6qcoo
mrYLMgpFUq9ldV7WWRSOrRV183+My4+LQIG6TsawsPsiPigmhbnjBnVAHgtxG/QMux0o+dWuXq9Y
Wt7WhByd6mxNl9MI1h4tjTDrpXE5bWPpNwPe1DerZrzFtZ3TZtJKbhANZZOxMpz5/5NXH6lJgNa/
wzgXLBFWLf9EXbeNB84haA/+iib9r1gnj0zA7PO9yP5q4ZRgqGGgn5SsUOz0Ru/SnRM3cm+1kHuI
vBGm8eBWxbLCRFBInj7AfBHCYeXZwMmIr028A7ZY+gflm21pED6WLvod6AKkydctMP/DfGEF0Hlq
uMaWk0G+mXo7wDng1OfCm13uAuOR+hqfqqT4WHAVZtLRaT0tzxck+D93tlUCoRVlSM8BGJlEJwdi
K0n1c0T5ZTMwrIH7glDhs9mjgbs8xiYxtaYbE9h6feVsw+eS7dokGYfVpyDImRbuWAbUpQgJUObt
KSBGMtbwJTb6W5eulCnGOhcKHNGKEywhINAJGjeZIDVn3RmJViL0cj1/gv/rit9g1bzYRRQ4qVJw
299jaMwBW2wPBIbXIPZdUfNDJvhPIUpL9zmmmz2V2KxEqrFUCsM/vuoZjW9vw1IBb/MYfawM+X4g
trFfEpFevWfHXlfRQYJUzgFkAbkiCD13et/yaH606KowfoLcQ0YDFBX6/aWKWW2WKbePa/9IIsO6
TafipbSWY/KhZBpys5ktY8HVW/abcTLgeZLakAomTX2jIB+Wu8eWBgjvo3wRNmCiWtajSBMlCLIs
28BmOrsGwN5IGGQ+6KCC/eXpMbIShqt96xnZa7ax8O5/j7lP1UxINomVuWysF7s1s+yPIhDqjVY/
MBiDz2qvyu1gRUo/wrhrQvD0SaKbnb2RjUvh0X++lvxiayGsj6Ujul3TuE7VclRVMgPgALfptNLl
kOL49ygeORdi9Mr4l6Wn1gZmrRaFlVRejD2R7yHKFJ7rxyz9e6AA56WLKz/tHbhq1I2ujmLMDj8+
Ijt5nwo/5LIfHMYV8VqKFl61e1PaYmGJyB3x9p0MQD6nh1i2iYsFgIfOCsQ4s9hLudO2KR2Y6cHk
ISSkYPvMZhL7/5A7nA2o461GLFmZr4ERsGKHlFo0+d2BbPDH/zfYPIIvCa84rgYfOEYBxcXUfXmq
cYqGlsuBwDmZQLpuwlbeO6kkUJmGCttyyw+6XIFU1puTl9GDsxO3zuHzvLCQC3bsmXQyPx4gYBYc
qXa5utcdnRxACmI2l4eb86SFtPfjf1fQbNgf2cHkz9rKeUZlT79XhHa4mjEHpHj9tH7kRECK7SpH
d+1uLBatirCAESKETbUP6Ofxt3iUlbN53MmxrULEPUCPBwultGxBgeL4lBp9+ZKJRtl1C6W5xi2e
uxWRKdvxy19fE6XP/DGGQaF85quR0ITNaw+Jw2aeAWysGpLOXl7sKRzW9ESRMzROhuXhSN29qIl1
vq/g7CPTq4FcV0jhkD0PTvAxjITBUfhLxk57YYSSu4qCtQH7JlZZIyxAkkUG1qMKD0MI17OvgF61
XvgsDzkQDypQK9f1m+q9HpC5M7jrOWfh6J8svi90d2UpBmJwWd9RDjFyJzzlIt9Obag3Etd74u+b
DmL8S1L0sCNYnBLvJPRmwF3ahg58OJosofaPE5KO30X2OkMXe5Ow5DMV4fhUmyytCma2GLUe2HAf
uuTs/NBVlgPdhkQqkZdjwJEFLp9LADl7gMCptvaHPyl853vqcUbY6NPBEOJmADNLVJTRY+e1PFzL
dg7ZGbFLFppYk9f/vZtLsb03XjUsDyVOM/RNuQjwInxZQ/NvEsjOAEQB98Nj83/sXyIe/wDyx0cP
en86zJRhx+xcSQcc/a24vqvGuLlUhRVCwgSA9Zz/2O3L/Tq2iPYKSXwfAGMRtsfx7cavu91siCMX
1A6pMBYgAHUXFXU0Tv2EWH+W9DKxKT0cpjjMqCMjG8PeBqjNoQ2xe3L3Q96o49tV5+j7R5K8wAG4
/vjxAx1Ze2hKt4i9hWSiYGI4yPFPRhvPOpbO31sPcRlCwKdrYZDXwHO98GfjndgogmKWKi0byamM
DkJSs6F7dlMURVtZTtDyPdWI9jD/dwSBRn7TKS4VC2xYH8z4rBGdBHW75/9Y+ovTRTxITr/TcUFy
irYIB8vyvKjvUAM9xemmTc8ztE1DbcRYBLMFo59iChMvGFr1QJD6y+mEG6b7yyqeZWo1OAi3c9lp
5t48haHUTprs0AdU1GnOeVjVDoxGyzmOd6UNwR4TANr+2Ij1lFgqc2T5jEQaEwTbbFS85lPm4VPl
5rtu6W8WTFwW9DgW2HI27Uvl6q9jx/ktCJR44Q/b5qx40+dbruyAz+lE/yNvr6Tgv3g3MxVJsTP1
/MxeivKQCDGY623E/JrMoWlwXLJQTfi6SpLrY2RQ2Ovr3E97IaP6ElTyHXC2isT+eo9JkIahtXyI
FcliK23ySzYXdx0c14v23jh1xbRns1T1KhBDUSSgMoBtJeNESgTxP/5Xze79HixVkCTv8Xl7Hoxk
1fYAoEKge/7ovaxU0mjJzCz2YmLhbka98P2LSU6KGDvMb5HZpBp2YZATDYlEot7QGSZeAdQuFEJq
m9eL0uwPNEpwmtna95wF7FRGL1slcbPOIwOnyrVkIRSHAS1zbdXxgOnKcMZLrBtCQQmdEkr2P8yd
pCJXGRM/QfcWT8WeWmE76KCWqLJskbEhFyCoRr6ZPw7J46CDT1nrj0/UDKsp2S/sUZWz/ulyZUme
6pjvaDOrWGz5bEL9M43XPl5xD7jwTOM7Ipzl1Q1TaQt+bxylNnai58Kf2uDrV5S9TgXYc9h/pgsL
b22lkoMKA0oaaiNn5jdH6hfdrKrVYPRqoYyibrtUnYGdIMRja1iZuDqgSKdksbPq7HCaIg6UfTo3
wxEWzmqiWJFCPslHvSmiQ2utW6ELqYUEM7D7BT3b9XY6f0WchDyQyxrJnbFgoeESEs/soaftu/8S
IY89SGrTj16v913XVf35IFhRwu3cphn2Ju5yAv+XbniCjg/jA0OAksbn8dbu9ZiQQQzXVMPsH5py
OTUQyZOeDyWFKQSegNesSwcxUq/wJgWKHP2yYz6Wm6wdQkVKMjJBAd5THUsKgctNtwsLiQOoOS9U
/ImnGDsqsHrvE/GZxZiW0zRoSM8ETJ/xV4VKZz+VauPbtFAdzHzhVKT/JGe/9cRaVAZJ28iTwdOm
aJsnLnW5LFfCX5Lg3ugjYPBSXgjSywpjTixv01tXcbKjogxbARk9BWHpA9ncsVOg+tJqiaFYwCrZ
E3x5WniXyin7QU5DwJYfnqEtUwrmCf9oCZS8JnLidSVoUws7Hi7L0XShtve6EmibSenQx+qR48iH
QhGf+EOzaTFFTkCXRJB7H78Wig2GXoJU+DoQMgBrrXb36iDrBUHAbOOC5fOIF0eSJ6rjbxV8m14O
VMd//YJQ9J7RCDUZjxx3R7lq1MH815+1ecLWEcLfvYmEnrLbQHJcWxKEcj1XqytHU/TI4mOg6fdx
mWoB23fdqXD/YYSx+WW5F35xqVa6SJV5srIZXGHD+B3HJ17Quu5id2OtMmaD0oCU177IFGizke6S
YZypUbC3a/NbncWmEPEBaxssQtEU9YnkPAXY4lJ5flJbWfn6MEu+B/OiA2nAn1MDDawZZCB8yiTx
kNWlQ1/pVLhMlLw/toKZBMTm7zzMluVQ3RWg507+dhZb5/9NGND5qaHSYuKvS0b76GUCEBdYnav0
ZqBGhGgyW3G214cYKI72++91MUxAF5BUDVg0TE7l4kc6hi9Yq8Ci1mNr3i4h9pR7jVZnsjLUee+m
q0GnIuPDG22RdLBNnEj4vf0ZVbCS6iuWaYrBuK2uV6H+nYB+fbjUfRUaIwATxC8XtAFL9TNICoK3
hGyB8TMNYqnu8bSj65JJZxqjSUDdKB2xeKmlG3GaVzSjTSXM0qAA+nzAM+6pT6KCUejNiblHemzV
W5IFp1lqZ4jrUL4UpjFkAV9bAWKMe8Esqld43dm77mjvDIR4EUECMqanT7c4iKFBcmrqsw/L4oyR
qmenMElbU1OdpwfK3UvrITrqRa+HEf7mGQ1vJ3MHCVgUxEqkK4kjeLMV3NYD+RWq+AQ79p6pIVVT
2rn1raH0jDrhhb4mYePa1eHV5Otctf35/7woaTBaXsgPYxuTPkW6ihT5AvdGCLPYIwyxejeEd+c3
jJkHHBZYlyx1bD0W4SKk0SGMgA6XgRLtaAeKo/9Yn8LBwb3XGyeQaCDAbASZLZTBCZA+NqaQxv/E
op+zdbYr1b0DPwNLCJXqZ+30uQkQjbka+TzIF+/2o1g+nV0ugxiJ1IzaFiUYJEj0Rc/f2bcr7ZMi
/NNY0QHNJAUlaEHuC1b5hzMmdZIvTbxe4ouPddOnQLKesaGya/xYWXbWwPJ45ucOdsaOekudPdKt
1Zny5q16EtmkQ8XLxPnhb3M1JkyC7xjxrPd0+DpZKkBHClQQb5jUUYLzEpqAG0tqq/48ZyX58gjq
Ma7t/mbTdWPy8HuMDqux1qBYeeES1V/EXrfyRyIdX3PCfMGFznC/yJktkgb03PAYdSQSDdY51Qof
dz3Lo5pgYx5dLWwAsyhn53qtaoBdd2BDUcORm/pd3xyMmOj84SSHJTsrcgLs1XKuBZwPdz25cgSq
tv0+HzpYZV9pSS97YDFG2eJw0TS1bfaK76DFZB2vgMGJMDSswb7EAm5O0MIfOY8Co4eVhfJqUuae
pj7A7pcJqgh5/hEGSNCSwvzZlZeKpOFy1Sn1hR7U14bdsNXhlrr+NNKuozGb60xN5aDgJcDAfVBy
6Mw87Hw4hrdumvL5lVyuQNLzUzbTKDzUVHVBTcsRw/EYhQE9wdlpa9D5C48uksr39QyRNqcsZsWW
M5XUaYwwf2/eHXT42+GcjvO6345uB80WPh76UyWBn/3uqRuseDFe71De8Hbuo7oSQ9Bnw9bNX9CS
cFzC3o5ARBJ/hD8bTSKZRB4sa90zP8lf2NhSuH3wk9bY057LXLWedS5TCBeaGenzCS9QS6fjEr/D
v/z1g0bZKqr8OhumayN6NJ4ole6CgrLHcasH4Sueif7k913nF09uDWzdbZNTAj0ZAjfFPeOWnY/c
ob39wPpzoLuJ/k8ndB+RHYeDgQO0KXoIfatchcHzVr9tkgmVkFT/VFBAe67Dec8NakwB6gsOIeQZ
nrH8Mth7hcSOLKKScMgfkMW+KJn+xLYatYY4Ugs91TLmI7H9q5ISXYohaCf3DrBasarexUTbwPaC
43pf2Hu7MHJX2v3ywHEkauysBv3x20ivI0pcqvszsigL7WUB96iuJMJr4Ihg4R2vBTdehPkvhpvT
X80lh0/MPHZ0L9QCeMOtrrP5SAnKD7W7QedvIRpt2trQA98aW0msHIEy3XwlqrXFgFygDabwFeDr
CY0vaIbR/2/lViUlHs89fC9e5jssmQaS0BYj0XEa2hqhs5oec25sMc8bxhmj9s68XQaaCRpT8T6C
BEP8PNDK0EXh9qYxkvRhWzXYuFzOgHCwj9jnaDS3hOhmoDzzxTZYtIHeU2DNpJFk9z4YEWMFNyeV
bqNvn65QBhJeTpjhhIILOXgk1BhGnCj6Mzq2d9e1BhYYYIqfU06Pe/p9TI5Fg9otFtNb/ybtRN9N
AECP7uSgADOIJ7Th2Aw2kbFZHB34yJyLVbe6cwM7WOfTPh2fSVRhL+0LCLn1ZD9qGpAbuP3SIBza
qQ/0ZiKPwClWh80tC9UPuisDEPngUfb3sER8/ZcPgqh1qHFGH3H67htXejJV4120lOTCKUSljeYL
vtvUkZA1MsKcllUfnUht8MEeyXnXtm0kAp8JMaRtzg1YykN4gC++slE/RFE2aOYcKgefhuUtfUXp
nP2TNjPq3SkOmporPfNE3yQZogiq2Hx8UTgoNxcpKKLLFLG6S7hqh/U8Yer84w3tx/oPrIaGFwyr
93psVYHk+eJhwKufdKyDMg7hAiUtYqOAF96LDGi+QRIn102QBureEoG+zSyO8amuyZ93xJAaMVlG
NspOA3krCpS9mhmYu6A/7HyzQ2tZgkpsNF/3OxEqpwNLvLu72KQJvT6jfFqaUGio7bJ7kCWVhfTM
D8yxG5aXpc7io+5L/v0JEwm4OoxxCHNHsk7pHJe0oeGSWTvtfJXvzBaw3/6xtbbRpNLNKySKUkNH
psqnO4rs8cS5YNggdgbP5jLhlbKXAlAXsat2lj5PFpJs3Jvnqa3x6r21U7Ano0T99Ruqy9JP8KGf
SbbHxqoqiY0vboKKqziawxkD4wJKE3U0NLBMt/YxDLySHb+MnwsagxuhJaRV3MeNTTqxsZB8k+nr
VU9N5odxY7u5fhKE9bBaFYYlGEOwsUUUeV7q2Fp3xcXrFm+5Li0dY/vg68ieFsb8UigJWEixaZEp
EJJLoGfVLFcRat4Bge3mhnLkhy5kcpLlgFXR+ZJ+4RawMSb/t747YPopC8i/8N9jGwPi7vyrgsQY
ySUgVpKwPX/Up2E2NG2exd7HJ7PIxwD5NunFSAtxeQbHWaFMpevP/VKM/WOaRsJjRPiifE+LFtvI
qYmjGmPOhwOSKhuigGt0WaQihtnbrvhnDyXYNJ+B/J2c7S8EOdvl0p8u9M7qLYtN5poBDXm994ay
QRN72jX9pIdnmACJX6rMFmSy83v9VLT2XwKW+yhUWSUX2OMlTsJD4vTmpAGYw+e2APyLCH6eojLx
YvXWjsLSG31xoNgeVy8S5I/PFNO5E+ohxGMHfcagot/h33xPKrecVqpHuZCuxPGYu+1T0FrVfcN2
VZkFMoWjQesA2toMLkm0mhhMVqdJYZhpKp4bAJVwAPY9mY4DSc/GDM2RhN/Oat2uv6qINUSO8twQ
1lwNKuaafWPGnJnZxE56JAGWOdLkxPYACwnMacKTgfvsCprxxm/5L0ilWYtOA5NWoaGUE0diQB2B
O6DEuHdEb3p0nSzgveILAEYfHCGIaWrynOmSrxTTuupqTs1t4s0DkwNlT9m+MvelGFf5tRdGmV44
TY2oChLQGURYGgHesRtgXKNxszlE+s+s0vZROKAHHTkc8fnsIIsyElcOC5LGFq4Ll5XqoftXw12L
VqbyVkrXnrh3JO4n/NewV/5jUMWZblknawbdPewKjUtKPPM8bctWVRlJFjpPdIzilKwbLGli5HBU
kqVqaegVaNubqgoD/jXCzpZe8z+UUF+KlVD5KOYyEiUwhCRCR5tatxVKKzvr5Wna/nzWOylfhe3G
9YH9hH1OEvIeVDD9UQ2UlERjjFuGWEpDjqFb1gEseevHLGtfKpBlXq4o4iRQfUVpvWFsi0vCaa/z
lR5rFk8mcwW3ZRNJq2YL3hlHGoEWuiPbPatfYRzlah+ql8kdKT2T8MmyAy0EXP3d5ogWvf+YG+Pb
CHhA3KN20nHKCrqRBldssOS643g8GRT7Zq3KZK1GXgT+4txsyYYtjCBPmu1fL/yDW0rKH4lATNHS
Cqq9RtHtkXE0L00E9rLIy2wUcswr10hRGCzW6/Es1DOWbMPBeXV+8hXqWwDOvcq8UCQELk+HOsS5
U1apJmqwTF2brhh7KqKjunT3ZNfLzgkr7NToBA/0i6qsDrJO5HYUym4jd5LSBaYdAmK5AUXCSJW0
VwaRHjw8RiT/eK3pdG9AU00jZOjhuC6TchkGGkMfEUB3cwIT+UT2dofFGrdWS0a6MfeZOLXph02O
aVbcvr3hWCTAFdEYHvITfpSq9AwdVvkuMvApj+zIoQRbEbQQ/sZceD3okCx1j+BC77c1B9AZ81Ti
2G/k7omjYI+/omZDOFC4wrXWX7VZTq+8mD5o0nBv1OBRYTJEGxG/YSu6f6tpe8kYbz+B03EHrC5i
hs4jxThO+SSZ3pOqSksDr4SRu3A6Uh6gZ8dL58ZWRXjz2/+Y16eOTxqgsMgbjcW82vJXKYkPFgOz
v7ZUAboiTtoMD9AppUI+vw15AClxwOVKPB5M6xqpWGGkmv5FmDqxzFgsBPtvOTMAQHCIxuz4cIhc
ZpECW8erPj4P1h+8TgG8JDzRo4R25rbwq26Ny/AbW6xFUgcWRm8o0eyaz7Wy4DWz3iiyCxUcei4q
H7207MSucZERyNz+dErsu9z8ULh8/qa6Nvtu70Bokwdc29HJ6KIBLVExkq+YaXfJuSKk4bkfRj/P
NVOuF3EPhcknpEwvQl5ceGUpKNJEOjKbu6UqlzKnd3kcG7oJBZIU7k9nzeAULxYjjyvNOiZB9xYh
Ba+LM2L5TLjCLKbVRrUtb2Olp3zxkNms+5qFfgh8mgDirHMoV/WvBvuDgOxrWg90GYKRMhOwr+L0
wzDV8Ur842mSrg9SGpMW4hBDVG2W7xCYpnaMHoI0AOpoEpUsVIs3ZHFavC3uZ6OattPlXSCBUu1o
9Pibua7HZpUGeh/0IR6TkcOaAmsSva5+h5xt/2GSSSAA1KOCqX3b5JZA8vNAr5ZFwKqv/k1qOl8r
GICW6Kksf8bEXn99FmPtUNpYyNskFXnP0649LbytXqTdyrpzH2znsFtU2im43fAer3GkAnRG8v3G
8cGggLUDKW/CWP4VkU38Dj4nPto6g2MxpqwDV4vR3ElC0ziNrZiIokeRpooeeWYfvgCFg/J5HKme
CVZP1syOrO0FPg+UoGMK85dKvmjBz3it+9pNGhI4OJiXS13uu1hGSP/lQP7Dr/HR8LuE01+Lztng
Ob6UY4wRBvW8QT06LS3R8T2RYC9DgibQL0KHLELp6cSBBf1r7dZKrDtmAv8Bj/pRuzqexCK1CEyc
rkcPdCLPjzlfFzujSYxRq1zjWHKMslFHw5JgbXYACyVC6uCnbQOQUXqiqUC05NKlsFGUC/r9LYOV
qkz8QRqiMsKtf3+iWGhHSlfGNX+H9/QP9MUBXhJ5StUSUdgK4ZwNgzhMR7qIp9wOlLqKCUnAsNbS
Feh9oz2Ed9YpSSSRPaD2U7+kziXprU7SXCVubBUBTFlgUvDdoEvmhQ+n56LtZiJSm1BXgGhA0z36
lsrqz1KafVqYHs6T0CfRq+QtqakfYAsdIQXPcU5pxIhqfDVZ7gPmuUPB7lLcQVPSIu6xMCWPn4gt
Ht7WyDQ37qV7ilWeIQ7JBOhyQd0rNx4dMJRrEhHiCrlojtcPREXL/hYtjxmTojrGmvda5z6xmFIC
r4Zb3OqAqiQZPzWIfXKNCQIQfxFcbVmvRgqpEOW5PVqNEXGMjDxvOKKH1XuTgA6/zvikDurrmnBw
gaD1Z7LELU/iKOszIcVs4G9RowRVPDWsXvmscE/R0xM1WaKgUqVOjd/2yvDZh/5Y9515c3XeL6rC
SGlSfYpx2tMGJMIDPsXNNnYj3fGsY71cjHDDiaU+vMLdKKXwcpavtD19QZZAQsvE0PDSjbZMwX3X
DJax9kXSQk/6P2U1V3P8MpM3S9HH3vgmfwGf4tM6YUL976xg2XlSeZVo2xDM0ux903dNzImfIkP+
Md7tShi9+8zWR/2Dc2TRghgas66OAgfHxY53uScSN4epkJafPAVzMToFd2jHorwXq4a9x64pYWKr
lf9UxZFUohAmGH/pX9IqcrtxuGD32BILoQT6GcwBsEzs/WqGbW6YTIIN6V3wvswoJitfT8GcpqHT
AyRoD2H8UBpIOqcdIy6mja4jn/rBOW4pbLSYWosNjp4gTwRLfMnWgVXPCJ6TnDpOj3O1uan8Wl5h
8eoj75LC1YTiWlZJcx6yw/AwlNuNbKirHG+BXfbLkP0eHD/sEQGxcflJfOYLuUyyv5XIkMXP3obk
c+RtmMcpbAAuBfHDIEUL4bTSAJgUXlmGCH6RBIG8/JlcU66QVNCyXe9aRUJcSmATg1BHS9OpT1dE
93GQj/R6LCQym5ea+iBp9TyXy0VUR++ICcVjaS9MFKCZT0KBEtZEuEl66zZ1nSYEOts+2h1BxtND
RUDOWiks5H9Do+Di43/leOQHXSVvBX7zp0eYQY157YeUBzIE4UVNQ9EPTX52JPoFXHkIKY79Sxyi
7INqPchEfHOqvW/XEEX3FxH5fUQKFLNcmq/l2rp6EU17AklkKMZy4rzP2nHRz44tBCwEzOBcbjJs
Gs/8uKck7r8gEj2lUj7HKgyPqZjmEWfUp3GcYApTqsIdZTIk+dIY/d2x4sH4sw0SBgTi5uwrrvlK
wRxKjU5tKgowXIsSL9CxApra+5w6ZUFKnh5Y4BQscTU4cBZyfiH0pyAG1XXMMFjRBm5uRHvIk18y
gPjoP+3AJHQDwM9lS7L7dO37G3Rc+MLX+WZOOmEjzSke4Lh1Jlcmzr6LWkaF8EncnId44Bnas2q2
o1TpxupnQeqlU5j8vhHRzLjthNpv2MmdmO7rnD/QUbJRC7x+4CzDTA60ma48+uzbkWblAlv7yumf
HaIwRGtBKtwApADCalkgAfFu6MzvJS7gqswMnQHS9BZdqV8Hlo4pU8THQEWO2A/f9iBwbmx10Q/R
lg6GYeoHDesLF2ZKiUPe/8qkeRMJ7jjwa5FkY6swXAgGgTRTTDVFXm7a8xdevyV5GzuYk0D47cNl
g2EwfgYCZQRpGQ2tUHaNxlft1oe7kh/PYdv7suIslo0PqYakCNH2QfI4/kzUItGs/wTzoFVzOXDK
AhS0Ajao7W4NXwqu1AZgxfiqXXG3Hlvy0mzBH5zeZ6dpSFbPiQIlwWCfZg9yUFlcIqzP8DdmosSb
/4/Fnj1MRe3F33YvSdsJvGsQOEHvw5EJ5MrSSMWTbD9r7UkBGfLpbb27BcEAOkwgePiFf67YPMAq
OlHG4A2UlCuvHH6YflCBpcQiHgMP1GuGR2GsD5gQPofO/rio59MJQvRK3aPQg6Ru2fihqBj7Lz9v
kMwSqSrx+I7FPdgSHLVH7jS+6d7a5FjRSuHOsb2c0gziy7fkLPv7fC1RBL1dD18v1WtXVzQTDFKj
35dIUYyHhziwosQCvmwmvjskVJvMnQaycADfia2N17f2SyIwMqjf/gEByGr890BDVah6BUx7ivpb
151TtGoFH3Ip9tNTX6ggpaz7bSusVNsbqMM6NtHwDr/AbDit0Rh0gJnOIleCor0Vi8U2OHfc/Tm5
JtjdMUvHZMpny4cp8LRJ+MFrOblm9QOLEdUZssqHUEDnoqwYbLqnCe/xYPd8FxJkqL7nukDLJx0B
jTFxoJDuksgbJtynj2ShTsNqP6kZSOsQRMQPHECZU51moHmHmbFyPE2o08RrDUaJmkJC8DIvIamn
iU+TtLOWMarAMeZQbBLjCP45MnHju/hcTkwDD0mFv+iBKn5M2/vkWX1Euawd8FzrohfqHQzkBsGn
ThJVadz1LOsg1AegIcuxnIU768i3EKyfjTfJiRy1aFlp0F+vZlsZcyKdEZH3uwg0Fz6WflleqArT
jb5lOAvD2fbrKTeWlp69DRJprH09YIZc57dLIr0Hk1MT++K6ePnpRyfzBP4viKukPqrboyVI7AY8
9g5PoVB3cU3njou1DaD+m8uZzUh6xeJKcqmctn4O86buunKHP0cawoeQNIXtzxAyF2LFiBcibnAa
0SGSUdgH4CS3jNZOrurcrQJ4t5QlTYp/lhNdlinr8df2r0FFRiw5fZnJTb3fEuK3287OUHO0R2lw
9yldxHYsLgDfnht6vX3RnPQGp5mzDAM/pdOBydIzHhVspz/O0Vx6i8u0u6FdEZpGHPxjJFU8dDCi
vwbWWeqebeR05IHsc7wiHYczgcRG87YMx3OpUAVc9zoRJmrocp4QWn82wnuZqNbEuLC5hUVIr6EX
ZJSoolN0X7RzUQYXWyKokwuCMQ/6CXiMLQNuK5UJMpAhj60FI8HsesQaakhIVgR98Cdp+o3annLN
A8l9iWB6mOo/5W5QMTWJbqYrjxyDz+U0JeI3xsfUDRujIuTpwLRPGBhyHgxCnQaVNsM9CqZJfwvM
DbZ5hCSW0X7Lfwe7wXh0Tv1X+9kj1tZWGwu068O97JbGHdcu7hHMUCzb7C0q9XDr2u1CoDWFLKOT
FUKTrmOheVFeqfZGYjtGj/wOzPTe6gijaffum8KwEucR1WARVzaBj67JaJ1f62Xp7u4tbJIs8BKp
VH40MK3ZT5hZ4TqjHs7stkN6z6zd4vFiKe9+ZxHS0U91NJFznWPerHr6WOHnR5BH8PofcTu3KkrB
Cnvo0J25AR9rkuC5czerZ4YXh9xRnweryrnfIPgOwWvQoLu82WJ2eqYOXY4bb4vjN9LaPp7MZNcq
3w8osdarzTR6LHbOI4ey8nu1QxzBVnXY7N8qZWKEQ9Fm8ihYH8i4l5T93oPG+beppADldfgkHl9A
yYSTmrrStWjDMRUNGwi9LTgGHJksTGIPYOec4WNEccE6pbluVI4rP+SF4cLIa0Rp0Kl18q8uW3j4
w5oSJjZaUqrrwyuC4rS9BwzkeBeFkH5b2iEwsypvUE3bFNRmPGb77GzxKI+zu3FXB8ec6rWjUssz
heAOoZVCRzewEYo7dYMVdw1NBb3GPrUzy4umMJmiA6YSomxdJnc8HscxZAQONzzlnms1iUR6VRMW
v6q2usw4Ht9dI2i6h3ChBvH8PKUky/7HUC/jPRGHJ/GZ37ICQ64Sly3kwB3xkbIIuxbPcR1VsRyz
ZbK/ad9t++U/23Ay0Mu9qljFvKEROgabP5sFLcfY3ZMYIJ/Lu+3Lh0T4viSuSAh099V6R97WZpGO
Z77MggumOSOsrak7N2ByFsatPKCUD/58uw8hHJjREP4mQyFafpRL1gKDwdr0BlBGsgKWG3fk8fnB
SryAJwpMdtBxzooWoH+FcXrjeVQ9vV3GhNiXkUwEsI+1wgCIBu4GYA7mz+Czz/Og+Tqc50aHiz+f
y09KBmx2wV3JgWJ1eraY9ZXwZklIGMkNXWypRGFcA1BicMYuRb8sK9hr0sMrxiMf5M16fq0lDoJj
tAe8jXte+ICv+uQ4YMfpKJOEbKlNf2lsSOpQlD+/3zT4yVRb69yz5xwjtoBc9DdNfE8Zy+4kC4YB
jwHJdqe4NWc4SOTfMnsDBSTRbvU/e07QbIrd0tIc2QhaWlMOxa7jOt+0qEkhjtMdnkBWF32gQPVS
uQ+/6mn3EAOovdQlmQWNOTUIOePDLZLV9otlQJ6jX1PCRKJiakLa1FwVU9f1L512Qo8wsUroqurV
Bzp5al3emSZk2EDFayYvIc/6jKehJu9jPCooNfi3cZhdptC4VL218sfsLCVGLLJQoOCNYD0eqarP
Q/ycibceiiT6+V8TwwS8t8jb5wZOSlgBlH+ZmmJmi0PP3WPUUvSRErSZmKL2Q+2TECqC4sjPCqJE
71ewpK0IpbtgPxEjqytghS9SzmLtwE88Wy61O69XVMoRvvIXI2jjHfG+ujSnWcNLXVL4PLHLfhqx
5zGMAXCztB5Hhxgu5YOopDRSk+IELE1qXNRUGUlF5x1gj9TKfcbt3BKCwIknfsl9t/w4MeTiAmZe
++cxyLE6QGgtVI6BwadQIru9z3rxqzuU/KWX3yBffrH/TY2DTNAH13Kg0EO/a5deqVtgosMM7u24
xzsEQB7J1vVVA+4dkkU8IPgpV+6nJN0BeVjQSgY+pSknw9znkVnPMN0yFtrCIVw8uik9bznWbPRf
BXMa0DIVxw9F2o64oCJkzAsMBA9OI4sYg3PNGdMS9qWtp7FDQVzQEHAnBtYy/mZb6TemqjvtHAG6
DViMLS8yS46PuomFgd2nChh/6tZzK4P2Zeek2NKOOzmphNuRDmTzOfat0jg1bvog2QzaL0cfehrx
MCAzXSpa0TRwp8CzaQ1LUP6Ujq6ax4XlwVSzy8pxt2fmljyWoL5GdmqNdmD7mCYZHvTPDsDPDZuC
ZdFRW6/kNG4tK7e75xpKQegvJbu95WFyDEYbM6H7YeSALQo9rwLjeVNARID4VzoOevfBNYK+gqlD
sqH4zsnzvXacywxm/p6htnTUYeueTCSKO71j3qQvsN+zIKdqKy8OE1KLFu2+L58JcCIkpub0uESv
NDzje2rR4HKVK7mC91NFNSpDiRHiZ80FaLRPZpsxmwqsI1SmB6JiWcKa2WfvDrA/cWrjp+mroMEb
SNu8/cSOnCZaai9CXmjje+JDIKML/dgcwsfcOGjAiK1dGrIJEItFwFmQooOKaxJ4O1nqR5VWr2AF
szivuM8e+g12xBMl50CmmQJJyC9Y3lKtHJW290AEOhXzUUjTGuOnBh4bKWbT2pWkfc1Kb4mjmjxx
wgTw4P4cxkmiqPtQne4LHE09I3WUeN/plTpo/68gN0Zk1rbFEbChNT1DUbmIsMILvHw58AYVmg5R
z4QLaE3l0oiHkRc8QEoNeFVVHxlfc/Z8EQJohLAOnk5oeY7LWHUpMtiNXGD1960wpI85/PwNpNg9
jD1EL4OLkKAC+YuwBVo0D+GH7PR08Q5MfPeWz2f2EGMuV7tBiIK/eURza9u5xUqSe3nZIi39UH6D
IFcfAy2CKkxb+ZRGl5xqlepI09hA6MSYcyoWfBIG3fNaAbJ8CdC7A4GzlViwdBuwMwWmKCO0kjx3
epMrZ0MgM33fZe8Rf7FXERmcCvKUJ74WbfbGhIvzFCh9/fmSR1Ldv1VcWjUxp7z7f+AXaYyZA726
wt+q1OLy1XVu0tAcyr8atay2j386qdw5FGu7mEJMBcXVC8H4G88IpgUttxC/hctx3R/JHukN1yDN
XIaiHxIHlk/Xs9TGJeLjEHMqCwVZPfPM+MGJgCkam5EAan4zYqtIppRyQ04wF6XO+Y5bYnRkGm8S
Fwn7GDG3tqiXpsyd4T/DxlbHrGgsYKVgyJxHKQEDmQgBB6o4oJQ3wownggpXbE+ffCZJnK79PGh9
xFvGOVhR4RG9MHOrhlPz7s+K9JDd5W6xHfL+2dLgjAGFs28MSfXlGaMX7ykK4JfSgOH31wuBG4X5
QjkIdY3dxQL6RdjHzw6DBIwAQhxJv5Mt0WFTfGYNJMSdlmmDX5C2mIq5JFZi7HtJOtcBa3Mqlp/2
a6xp85TY6CJzrZhyBeCXzGRQhYlar4vsVjzbmsrDDSy9rct+TXlQuIfatSQym/GbUvSqJ7vC1buL
EA424KT59gC6/2AmchryFj10q+a8KsKXQBfqtX+KGFsMmd6+TruOdSW9t+Z4UASuEtVcmg1U9PiQ
tKpKEk9IIGNo51K43ZdPYu4BkGTAnk7EQzywDv7y+MZufwxpml9XtCDNZk2U3pZaKSX6TnFuxj7w
g8xEqp9YqKbPoB6kiQjqYwBitatB6oCHzgJG9Ga4G0wW2sLmssqMj4AhO9t2dNhDh0yFlIrIIl3z
SBwoUfO9Wc611gsW5+oBzAL1+ZledKg8PCzlmuM6hDYLC3aanlcY8bn3RRo5rVJmVfFIwj6fZVUU
ZalrLT5LsTDmh2M/ap5w+o1wASR7zwrnGQzj7F4n7tM7WaWZrKvl7O4S8U2CjMNjIViPH6wpfA3G
wHpM1VDtLElf3fCssNdq6tycp7abHlPRsUjUB2hq106MW/bJXZO6z0gr7m31GrukG4BAU36Iwsbf
RCN0ydysMMTV53mN/A6nSa8ODrAut8ZFoSSh/MyLekLNSm/qok9QdRpC/bWswftiwx7i+dRL7jQr
jDPVXmXp8jj8/+wmp5oCYWTIO5jROuZc51UfkGoQfZFE/K/3LBsk+4ldmTmrrISgQ0Cn1PucuuSt
w4+GxNJHVOh15a6+e2apkDQsY+uHJscF3nwC4EnqnF69V5SwNeq/YNcEc9Egs2cLynKU6w7KIj/w
P0JESOZMmgxSxiWjuYavnZ+OZBT1EnvV+ozun+hEvZZJKULiDkak2AcgAIHHMa3pgEYFvnLhYPRP
AntXWCikIJ8dXnjFfxHV50ak/nj4ed6AAJVr35VqphWXX9klVhV4dTLjhrE3BNUkrdbOMb0+3up/
LszakqAhx9EwhOzquXU9OTxrmx32hgLA0EmRiBul3DlribzzKIXGazhnYVITvn4mJntuL1Xu3cE+
Ly3vhSXPoSWwmoCBAlEhkFqdW7oS4SftDsN5PuGi5Tqp5JE/FuerbOO8D6wlNn+N/bcIhCU1kZFk
w26bAqtXQn/7ug1OaYdhjqG5/KTLzTD89skK1arTlX/raq3UfaDhpRtUZ/RRZSIxiHQW6uZyhD5L
tuuqo8W4deWoXKvMvaubDVB/JCcuO/bIZFfdLP2aGhuB0U08B+N48xZVXcwAbmLssJYFpkt3Wxus
wj1Mt8wDQ4EUxftQPHuTsos5c7X5b3HeLmuN/xAZRsqwgTTo5Yf1o70Kp2KYV4im7a9wHdrwDzBs
9BpDIoRTgfcs8nIAtoE3f4Gybz50oqc/OeMZjeLqmvWNwYNEn2XJZznqgXgDum37SLmmavuoZWmc
wiAKbYo06QHLc5Y7VpOCZba2nmXfCAAtDqj+HbO/hR9l38maP2HijOzPkpXYOxgSMG1xTrUUBsLk
yPfMYVre+1VGV4Z+QgW7EAt3HiAFiS3Az8Wtt4VbEiqm4giCh2KkESd3JBH0JsZ2xuqIJ5OyNZxz
m+pygPM3dVeQBp7+sAdkMblfsUYs8ZFEjUyIn8aZmMKHXsC6mshRp9EEyIty+hu0ZxkIX7NDvm8u
GCH1aBuXntTMZawJpSYcdvHN9z/6gtYFp7gAkVaaPz0wtSJEhviP7O37hR4mzEtesdE8CRU+Qp0r
TABArMQbHmeMhpKBkDm0UQM772rb3U7LZpCqg+bE/yotihuhfVCuv95c1Lk2VJEka4bLtf1mwWtm
etJwiuAklCUfn1SMghX4WGBcik8qaP0JAOe1DsUFmWohboIi4NE9qDjupo3ENl6V+WLa94+J4OzT
wbv3mevmex4jEzy0hCC5Xl+c7bueU61bPJ0Z5r3IGRyEPDS0LvuM9wTi8kmgRLTmrQnNTJXwxzfc
lzTAVEfocTQNx/pVku9rBn/2+xo/H3Agza34G0Cd7L9FJUGozis4uXg4E825Xlj1jmKMaglfxaQC
ycDm81S8MMiOmsas7QSB3mCT7goWsZhpIC53DTfkXKbnfiM5qu4HfYVwIMMVpLn8fT/fk7APhFKB
se6vRvfS4r9DaGDGnmsPGT2EtA63+i0jLNUnNpib1OJSY2bSTTr+BXobtP2WK7/96OgyDDbpR0l9
Y0HtComRN1EVVfGsU1hxSSEHyZKVIX+FKrVUAqL+OZkOFLHDVpqOWgHddcaAbIoybLpcvHTqHRlt
7CjmvEhlUr6nk9qLIsinsRs21JC0mRcY2xzGOx4r4XS0Bz43L9DKTDVvZuM0QQNLV0d8Dso4+3MK
czVl1xf3ZC6YpLp7J5Ghaf/2Djgv4m8jJXvHRf3stP7ILtq343LXhUQ5spUgVuQybn6XmFepm+w4
6r7mvVuWaO33GKnH0DYXa3pSf75lnEoddhsh97RJcdkFT3vh8lLv6aaSF3LJyZ1GucF7mqCr8np/
O7MkYL70DYPwKEVB0dP+DVCZ7KGyW2mDwN8eezHr3sP8fEn3gro7iuTs5sRMehR8QueG6uqREhL+
AtIwBmYxbcWm6EviL6Yz24oDZ991JvNOIeYmw1NMZKIAbz7R5cjE7fhJs+sjP4lLZqu/LwTXWtfC
pstPAceEwh0io+00ohstN/CWwgbECPU0Bmg5X1mkirs11BBb+VWxtqpAmcHOMb69tlLDa3aqKW60
p7D0wpG41d9lMshHpBrhPkOEhIxZJFNpr1FKmaQ7LVJtu5z02t0MIK2P1TRqqZiPcMH/TvFpaZEs
0Ruz1CAR5v5YM1pfYSW8PhyIwSvRckqBRuS3XrGG5vVb06/cPrHG4kNYuEGbr2ULa0coJSrJw1L/
u0OTTQiiGiVsXSAIv0DgicMG9cu2YwN7qAmLrZ9bXplLy0VwkwBgn+6/uQ8Q6xwjYQj94AIkqGbR
mNMj+9Yj+J1UyF/gNp3VUl/NfU5hbAG7txbPFBr9OGpLWB7NAjHdCiZ2wOOqjRLTaXdzOqLp2a7r
O+cqT9aw3C/dO3y5rzJL5Oe5iyHHaviwdOR6XoKD2rSUBy50PVIkmhCihym498zQBVGNmHkZ6P9+
uZtYS1C61X6MXnopiEYSXRe6qajgZeK4ulIYClrlypnAYXdJi3/en3IoncyzZHFljMbYkOAFb6cX
i4X9ogSkze89Hadetjng3HCmFwRa4C1LSCnt+FGGQhcngMyvjfjmdWsFGLdcb5XQxkj9MILfhXL8
N+cyzZOyqWhfGE2fxtVZnllyRTDuOvf7Ph0v84tcDtP1d1/ZxRVzJUjLyGRl6tHqCGkACnvFo1Qq
dXGzpXGEzL2lUq3Fe28Utba1XIAhAa7GuGC91vi9dIEuoG5fRZ8z2u3UV0+wbvnHzUTqmIXLPVbj
aJ09l3uVVIwbj4I52D3JrXHFNpv5+CrnpGJskA5Zhhsoyn5S/SXgiWHXApLP+oJJpp1z5pNPD1Yh
mlYTkCF0NKqqzcxBFolHywtq74inn2W9GEyRYrMvFO/VQAjDGB0DCOdVKXImJkVPtsv2gcCxJgGe
/0iolNcf6iJv5dDRFVb7yZ1F8KvJk2dIItJVyTSm0IuQl9bpkS6y6XhllQf53Imlp3NTVB7oaWmi
60bp087s+k/4AVHjFQXFLM24uizM0s+qHs1eADacsMWXOsT/Vbchg5gofBE1K8dM+jaw6cl5Ju/O
3HCZPjRuH7kEFZrlr2yQRUkwkqXlmnvMxT3sUwvRbllQSaz+iiNFHTD7XpJmBN+oszGZrW6CsGUZ
UCxw1WZbdmXCSQuxtZMfHXF2KhEvyWo+As3hHRmG/UmzMV8xGlldIBfDDkucMl9ZjZXy7Vm+cAwE
yyaHlNBXXb1Ov9Y4WoNJ08KTr8vq3rC9FNBTILPxyP4p/11Vvgi9wCyRORSeu/R3DT2BSUhTB+rt
xswXc21ozgY3qShyXtUOxkHR8WEhZE/9PpZpgH803ZHTeh/QRAdNTvktUU7eIHDHwrmZMJtgow1v
ole4YjP9e9CNyDHJ9Wge0J9Jt6sfwykmayoLovTgAC7OAztPdMHloOsWQXYKOMAcEkp6z8mhUcf0
thDL3WpM3IOFcfvWmRegbybuj8KH5Fd3xY0e4fL776UhAHuZS/VXi22sd9VC1Oh7fMcKXyTpCQSA
rxDJXmFe6bctPFeb3o/tcUNsJ8x96I20GMdLSHSEbgrYEkrblOoRZxToF6vKaaKv1dGsK1PW+bjh
CTb0rCy7HmGSJ9bgC1LyIv3BYPkBvRkAHyYEIzCbQgQHr+vYW9yw4I/vvkFycorT2JiiwTLY4sWp
Sur6gLaxtUVSTtyrqayXx0kWrAMHSdM62yVGztyeB5DPiC0B74X9rWSLV2m3t3y0dqzQ7OPtuYZE
e3Y0fhaWqHDNXU4jEhqX2OcAgwUQyf8GHHsBieswzmmYpzHvVeD6KavFG9lIrlkmLfT08TfZewBY
KJaJWxbXJJ9MWEQgnyoWitzDsAaVpE6Gnu9Y7JsoPi8U5eJ3K405mhG+MQVbyikP+7iFp67gi+Ok
NwhKRNnW3QmTBmKw0HCFlp9tyJqsD5YQil2ajAb0wGGUod3wClBRFqgU4lz852KOLzxjO8gASq9s
uu59iehuc6kCotsxGqy4hAO7SgvoDbMeGTRVKP7R7LipRplRhcT4gxQAXjowZWpDBSzpZGiNrmX/
CprySgQyrm0apvyamexK//WDUKLjgW9EBj7cTa5xzAt2D/oR6ErPHJ4VFA269+VH9wkuFkYeoOoP
tDBwZsEpJVFBd4cB9+YaYVD8od2QmjCwVVZqJYK3M41Z0xmIyba2BxC2zqbRugnCNaRpL6x5Zzy9
iMAJgSIRnfbejISnCc4d8dhMSKF0bMbWfYGkwnKaHi+afTSn8PhdESKhUq3yrj4Ip3evPDi/I0N8
CqMRUWSTuCdz3RWTkBpDlGHvhB2x+uA3tgw8E8uL4MpSrYZMcEP9QXlu1YZhdlnTT5gVaqQXxpFq
Ila+M2KBtQzSzOcoUxWxKpBIZOyV400IgY646MlcYYrn65zvu58sE4K7C5Gki8fWmVzX7G8L4If2
UZ+Jl7O/XROLvLYWmrRQ2q95wea/e5Z2BZVLfxiXLXBPRoI6mraFCftHESEeh44en0MIZEi0xU9Y
WZK9J1UzI9DuVd9K22p5V9VCB61TEeE+ix6yxJnKR3r+XsM7wEWRsVynrIOtcFFQzHjKw9dh8r8R
dxpxje5PigUbGxwV1CGr7YjQ50fsvGuAw6moXLik81zSvCe3Ii2BShmLzeSGCDoL23pP+6jo9OQ1
2AhyFvEc63AVhgz+wP6kX4NJA9nQCuVyGvTDBV/3CX9zM4GR1gCKPh1/yqWeZ87XAya/UxqDKaS3
bFQPd5qmxbSOyxU+s5/8USyleD9CY3ot60OqzJySNVY8BgNxbHbLpgoPHTIbPcXidiCjm7tGOuv8
3KZlDP5UtjbboLaCyX2fLK1pZByYPUlNxcWYP4HFjEAwCzZGC3D8rIgd0OsKPK2KTn+zFE31YIzA
HNkkVy8rDu61bhcevouKJ+p5IAe4B4/o/YrWkVZy8rI9b9vJ0CcFH6My53xOpkg7HXri4P1dSRA4
X6uoKv3XjcZFdOAsW2EVpvlC4ilbWsxAd4NyL9Unvwa3Ae+U8l1gPfKKQ6OPK3n2fshoA7+bZ+xJ
ERDA+6s51GUNVGkrUM6AV8y3IjLLMgCfKQgfxHmxgky+IPeVeL7n+EBwefG1MIxR/pCLKAwyW6TX
zDGed+cF09fDHhHUbccR4xQynkapiI31QmJX8bCPSw0DAzYiJuulbn8GSvY8OGj+EqCgOqEzS4dF
PUFUC11FQ2Lf8uxfj9ZypuFZ0WQj6O1pGgb+mrbY0zirUAjDNZeqT8y27Me60+RR4uwajlsq55K8
K/h1tHl3CSVOfPqJhW8f0+sjH1EB9fcItXCPUQ9OarTN+GuhVZ0/BgX2ARaxAjLkIR2qdGoR7tQa
j1A+wfgCycAcp9gEJYYCIpFiWRDvkxEweudzaC8IQeTt6wkItvOe8VFVHBcfBHNgofEZlr8uPHWf
sdE2OKh6sbJjz20KsOhhsW2CmJv6y8iIRew3Uy8Egd4uaO0HY8bXBJKW+eqjS+Qm7+Rk7985vdoU
yuh/kKh25JQlni+N8TbAFYLlU/nGA1ASqgdzmSCS84KN1jM15XYyuO21Zv4bfS4Cn3L6ItrTTwGz
qp1FueOiaPNP4IdxDiDPYipNUCMspJvgzqQVK8ha3Bi6Dsdh+abw3HPI+c4Hm1njHQPsqjvX2fSH
qPF4Ja4wygR5VW6SpurlmwmSsBYGGNpAZaR3ko3fBPwQ/KHjZf8n7FDUKRAPynV/bSCvsbjNu47d
WT91L+ME8i5PhGYJBfxBTxrOSFfMl5l7usqk0KqiUmBt+hjOHneDdxD2rVTN7vHFbC6za6v+CY12
UqXQvV2WqrG85HB27tNrhhn9ggUZZUkbBGJrLqKwkC638fb7qXlkR7NJJ+By66pDNrDEN0+3oYyy
vgHABmhs75JR9XJM8jJkvUlkV0PuPuKjij5EtCQacBCzP0Bg6aMm+I2FYVkXr9Pm/bFJ5d75QavE
kFB+Exxre4k0+I8Km7AagDZOBvLAKKX+0c6uloxwXnHYE1FNHKau7GdTNoel7y6zQeYWtMmgOHDq
9s3uNN/KAu7we9fuyFZnL18Gys0imkMYNuPiNGUL1AAJglkyAIGCt0Sdj8O7os6pfHQ66VF4kWfj
hxAYMrvSr342fVmTp/zJlgUawO6xdg3R2rtjVUlqJN4vouDnlU85h7oDDvT63BNrDSVkVuPzShrj
QSLvDPUWfBXP2FnEJMm8zPsuHGg3J2nXgnt/NsDwa56y7SBvWEvi3fUBqFjppdXWvYqhNR6pwQ+W
e8f2FET9l3L+MqN9tnaJgMV8HaUwBluWmPhg+Tn8TzqSuxP61WwHSn/lNiXY/xw83iH7l4fuRGHE
4vBvb92RrkREaxqyxAEHhFFXpvAf0zG1KB3uZolrfcdJ0HlvYa+TF3N9E4xl2GdkKDlD0zoPd1mQ
mR6bMVgq5j72p6ddRq6wO/dak4GoX5IAleB09RjTmAug7HA3rQb5nITC1wH4tvDiGgDjB6aNTKk3
LpWAxHLrfb0pFGYh/JQrZN043rYjYf8+zMmgbrJeMLV4XttF2GBQIekWBiZKjcSaAA0SRZjJbQqu
8j179I5i2tTMl2H40BxUrxId46iuBuz+YdbXHVJjE7vNKfs/0jclPasct22R01fzfrmDztoHkS3/
4EO0bkmBDyz8iZ2fxbypayEbCW88bcbLD4LvMJZkcg6Lmi1ttS2V51U1zO/K7ITFAdwnEn4itWBA
cNbhVPIgyR6yRlUoG4wpsmkHL1zk3mid3YggQovqvkUcS76mGEMnRWNAuYymvUjPmvvHmR4AXsLf
f62Rjhq2cDN1dClOJRLprgKdTFGv4ZlnqlMwOBPDdNX4GSArl+wmgpUFDCZ1SBbUzqtzSRqzu2mj
ySj0SDlajb2AK+cNIbzduhmrYHVt5puC1posyITR3jCiiBLqKXIJmcF4Itha3UeKu0eeTQY8Se2c
d/IKK2Bg7cJpHqHHQ3Yh0ioV4HX90Rl9kK66jTRmQW7jMvSjrsn+AK0yCIxDHf9PCj7QZq61kmUE
13n9U/mJYewNlk49+hx2ozJFxVxyJAofLLXtKJojcMh15uSkT5W1a6B+AvM3+wKCcpMU5thvsM/W
b/ug1wouf3UwGGI4NC6RHaaBVPcpmlFXkuhWNHdzh3BmUniBjEIqL3vey1rz9QC9jRb41ZdVcvFq
99DiJPukDslx+VFrF8ALfaTSnvwmgHsSkZiU5JZr5azGJY5Ku1B9iZgUtsAW4c1cG6sqFDX0rZYT
L0LGAhWBNMqAp+oD8jyovKeMWQ6WLU+7RR5saLo1ArMqSbn9ia34CG90XR2jNJ0MYno4IJ9p6z46
5Jvyw6TsV2O8OKNuQ5y9s09fGathjkam4wabSHTvk5qNUKwNzauplW1erKxOYP8IyyX6f9S6a96S
t5OctNhQW7oG1IiW3wEX+EjyHLe84QMAImt55f1Y4cN4USx2scNlWs/jgUiPDn135ze1v/p5vlvV
1GvQb7EWMiHJtmq116/8coANEYRUp8WBEkZKJNW6C7Ob8qk6R/B+dnh4nsNv8VYCLMTDTkIPObFB
X3WG6Jw/Vv3T8ylIo2kCxQh6Ju+bBKAtjR/jbPJg+GXVYOnWN7P5SDPOUss6jGmfJlDOYL2YPx+I
mD1VXgeACguemHsBjpAmjMGb1Sezy0j6gqVgitSpNPiCMvevsrcCWi+DpPLYI6wXasQTFao7QipF
Mi6Wj1SonjgmnqIWXJx147fRXLoGpN1RzGb9RFA3xhgJmvIHpsvg6MijYpSASpRBraoZiS1kzats
NrpHOlb6DBDNmQmGr7JNSEv33n2bESe0EPSrpszfLxPDLZo/MX5pySFnfKamwVDkCjr1cpxkxncx
hj9NVinaBKq2blOu1KkPtMzt+HWfax1DQYjFy1jOvcXYA1g6EDE5Lc9+BwVpligmH+Wjym051M+E
4wb+6dNer/RE1h9SXMdBaXSqPoNacBwAQ9GX0KsLBEfX2+LHkffqYyd+m9vrFjmW8D0wFYa0z3qR
PrubL9/dPj604wF3JoMuhkGbxF/qh34+2/dRhjZtOEEhLgtAiY07EonFTxGhaEraXIW9ZFjyvNjq
OvAOuH0qp7/aYrVO+COZhYzonRZLUlnz+VnGoEx8qKvSA/KamXuRTAyOSncOh74NBGblZBnUX6c1
YZeP/Z3l3DHEIMoMoXPUx+zp7qtoWa7PA3mToOmwY9WqS8HqWYucmPyASlAXwfvbdheWgiLWxHzB
dYfuNq0XRJNODuwsBJdzbEQMgN94Hf2psGcHOlIXCO2bWsik9a23IBpBrgmIBkdZEJ209UWXlL+h
NyBTcpszh3cz3rOPLNEcoxEsN0JnYep9Ezhxtd9kTIg793rMzIaCMBA9SRO5F3hWYVc0qsavaNNJ
yufVeRB+FNcUZZbvOdS7Qy96jkPwYRu44KCG//WwLr9l8lPRnAlaFeSwnLPtqtxURZAY4zjhgqHq
ZuhdFTEFmlXyXwKuz2fr6RDRpJJPqNDuT2vvNsbpwAobbkmRIDFOgHuZGm9HNrlK5qA+vP0oG7YF
qix8ZKjxgCzZM6rJ7p5cBmGEVRwiMA8Nt95QOlKvjg5pjbeMeV5qlnPqUmUG582CVGlkKS2nxLZM
ebowZbP0cTGPA7n8CVnRRanSLqOxMU+2OFqI7GuUHr4p8CA9J0otDQ40tD0z0zI8+sk9w9hwhOtF
Nh/5dIOFg0tOGHUGntTXP4luXSAi1pQeG6STyYIC5Z/i5VPPIhgMotE+7Abj6EHcuEaGZ0j2MdLD
9cyQUIwb1O9+TAdoE3Jmh+zzapG7dZRwokOkWyi1I3Z3NgnghR+xSZFJE/gHHVsaeBTBydN5fbgh
Jh+fK2FIwVARQcgV8iC8JMW+4zULhk78ckjF6sdTrrsFudBWdKyFuMGuvU8j5p0faxJDisogD+og
aqNRt55FWm5QkArn/DxZ2YrZe803tAiAn6pbzFbQ9B5M5QRKZmZEsQEy6c92QkY+sphpT73RpzLa
fBPS39vFPKfaNDVysHV5u8Sl6L3DpnMPAADh0p09tBksA1Dvu5SnuH6i0MNQPVH8XU2D0ZsIAgMG
p/O2vwnKKjE+6JoNB7gH1z3nXVOolCC3p6rjlNTAoO8AeMR4AirbSkmN06DE3AbXAguMGgO+xqJ4
5BELTld2B0kuoTdfffQWmruZ8Ks8VnlbJr1Y2DcZSlMUpxthRa7JX8MpsrIEqXyvomapyG9xjxqK
tAFeNrL1zfSuX26J+dp1EZWmCi/CjsWjOsiiEUMiEc1Vzd4+7ZhtdPiUAYuT3CkhgwOWGAFjAOrH
syOzq15TucovKiXpx+/RE8hfbyvNQ1CuyfjTfZQ2YrL4l9HS6kWMCplldSCjOJROAK1C9cldYKPw
0tAv0hvWknSDWIwSr1Zc4I+lXJUqdvt+utHzYAHGPiH3lBFxGtQSwIhkE6xvXtpoYJ4TO2VGefBf
hqihnKOGKGu4/K8QHgBNXUGOtgSKae6qcGp2zsLuTqD1P9MQ0qQJ18XElLKqqqLCZtL7YKKxohvi
AB29tVdlR3FsbV04VP7+/IGt/Ebwl9pQ1W1paTktZNVPQgrG9PEjfK29Ld8YvgWMDl/CnMfCebGv
GvpsbAhB1xq+IFt09b5X0cbwzEeKi31vmhbQv7IahQLCUiPlDM75aGiL8NnM1lW/BHPUwVuMc/hP
muLJ6OAl7ViLf3NYpJfZbNJUipv5K58OzX8fybCUvqvou0ynFTjEUZkSu2ku23eLHcVVDEXSLCIh
8jRm1Dk62Yj3mcTldtpLb+QXtKb3jh6uGBgsOGXewYtp0aVqu+F+WTBs6Oa68sbsO2bI7tDT/lNy
gDrHY5vZ7qPWugnHnoL802ddn1oG9/KHh5zhwFSdUB5gBgjPgHZdukEMz9LnaeTlZWLeG+i/C2+J
eMPxvRETlP0Me2RKJA54v3s+KhGH/XzQ1y8cAGF6sgeG1XkbL6ZaOX5OAHTzcAzg0zNP98UZIfMA
NvZq8Kksbc87VMy0COfDeMw1vDo3Xih6hAMZAJiHtlgNhRcTmzJenpamjk8xTm2gEU1uOEwXOrjN
9iyH0oet9LD8d1xfcALa60uPW9QKC6MFgvyWsU6nlgommYK0NAlisRKB05OyMH1lvOs41HOOOsDh
FivBRO4BXYPYyCGeV1gY1MVSkSl88DlRN4Fh/ykdc+dR67dfuTWO9gYtDFxTAChEtOK+4Nc3Wl9i
ozpVIREgPeNWuLDPkOOR0hFTwTvl71UJeLRLdxu/kwSgZX4I/SPYT5dsyoINxKHM5S6dlLlvyOJi
d6DOQfyerK0N1KQRtqgi6f5y/p5xgnt4HSGM2EfAPXjxCKt1pBVtdfTSfZMrTQbIVXChQ97qdANJ
qjApC2A1eebMsIZkt7+qGhhQnzvEjaOoJJBQZpMfKRZBLD6lXi6xWwD7Mw5OZig4ysO0AK5LFT7s
X8DxkNumoOqHbrOhZDf0DCuCoeQ1G8jSUACOJ8pkAaeiJ7ij4pg2MQn1ZCAL20NJLSGI0lV4gRAi
sRsM08ybKw8+OIM1q4QDAfmfXMHTF2+G1shJm9pLiS3akFjOTlyEqjQ895Lc5xkYFUBWAW6uBZOm
aU95Vg3Le5WGEgH29Uz29UNkpbwkXmLyryk+cApJndyH72ViBr57W2nZ20CyQb32CFbeehAYVg2S
zGfmhNQSbVqhJvLXBC6ThxEauwYAOwPGCt7BWjwitxbJIIiF8330e0D/HgAzFjVro6lBWFNynIO7
sKW1d639hk1LXE3K2r5lXnad1+idf3lVwlxj7kLtataKSeBBL155LacDv6sJIuTldrEu2bYY4At1
ZVVs4xeANcmEIhgN94hPoJ/ppP2JeY3qNiOUaeqDi1IqHiPy3Slh9y7zmlGz3zKk487CGc9vrMda
gjoypi9uFK0igFRyeqqiAii0yzHs6QtV1YC/mAweb8nVDEgLngv+cGG5NZFkUbh4a1xVajixPIAK
wscWiG7o7Jje8C/yG+EqthG+dUONQebkUjBmAKSqH8zbICyeRPyrp4vIsiVBHqmRrfgV/Rv2lISZ
ToQ5O6QxwxWyqP7dMRbnhsNBrpCCO3VtdvJ0cIFcqllrbZg0vlQ8pXRXswJMgLf3S+yt/ryx3tyA
EN0yvmddz528imDv/xNnNcklBZVTTFkf1TyPEkRl/2Mp+dPPnbAQ/du2SRF5di8sds4DBbuuBAwM
SmTqHenOaCh8nbL1RdjxvxbXgTVEy36EFiF0CB1p3DEQr2t2l8D/l1b+hjpFKhQ10WtrYj8kcDc1
soVbiVg7wt0WVQArmZcuJTTwoKkNZd/TYL3UKNtmk/L8DNsjFuTKv/5FMZstFTYHsgwfWFV94ETd
LMAqdsXcMDNH9YQ0Nx79STOvKLka5zwbO8IXAd9G1Xwf4a/N29Yn/7LT3Ocj8h/jX+spGxmFr0nr
6EdRDl/hH3pQR3hMg33wAxON/0oKVvNw5gljiTinoNodApeEJkQrv/hh2Erj4TL4CnddPdyXxgGL
oKrvcxoemLAbRMHlj6FMOquFTl2zEf+/Xtd+DxSEvRuiSWlqC42ISG8HpYDDXwoRiMr5S/rdMZHc
98Yo39Hny4XB5/S9W94FYpI5ePFTyaXubDFXhORkMUlcq0GyJMy5Doojscu+4smVS6HnjdbMi+Ih
n4v5CGkf9MGT7KAfiAlXlroCgmuyWN2/9LSZbiyIeG25D5qiZgu29mHcPX7GsFYhfaoSXZuKUWaj
P3x9y087trzultoZXUiSBJQ+D7Lh1DxXjehaWzcJkyyFKGh0DBb0YnRNiVOw1Nocr4FDdZDemop2
rKyRBnaeGtntP2Wm8yF3nPLSgwv0iP1VQNwJSXoAjHKDDPoE6U6E8duFiYqdTDTv8FUjzREq+8Tc
Trv7yivF2gLzMEFR9RwH9KSe2gblfMZR+Md9vbV84nlPulWJ6C3gWpB4wjxYBM89rMFrmMhhxoGJ
2SWz2Fxc9w9zZPWBwn0AWKEk6KLintnQqsR9g+OzZt1VrBFogtonOzAKD+eYpT2lhr2uAwHO5ER/
5x15KbUXIwYw0JJdTgnj5FmhOCM5MxPpUhEVDyzTom6p2gUXkZvGVXRIh2nrOvZNCvRTmbZfg62H
MEmStD913DPEyXeJkanHXrxxF1tt8/OW7OomP9Un+0zn/nzfovB5jmjROr96yPMvnHtgmg5AGVBW
x788Kkp5GgSuIIIWMWHMIbTg/cLWUNz9KT11bTvdk5gbbXl8hXtFiUPPSYVdtYpCKZzC5TfnvSXs
PZQeTkPUJjnmiSEusPsISFe67IHAJRj9l1rJA+qp4thN/363ziivtOpPtQcnoK15PaIiFZBphvAT
a2zE+FjdnQK0tIuhbZCIss8Sg0ObfpLQo6+K+JX4ywECQCVdezcRpcFGRapwaRM0qXPQcj99e+xS
hKUJFdlFfCQRlOkxHNnJufhgDc5b3EU2UTuLUaGHcJVd29yob1qyMq89Qfc7qhOhl9aL1pkM/Onj
Kev50JHIhVJEoHaFHUQEiRoy8hNnWghObA8O4X/TWl5a+2YaCtbwT853U9KoQRIyDXY11vySjCOY
PdYAvoj7xwW+C3/mKDaJXSQHEbGkLXKP5yxokwCgxOimCFBdEPDoQAzSKHnQ9w9rvXaA+W3xjH1r
jqKCQHN43HoUeIWKIxayZ78iHHc7QHN5wQftX4Uvw+t4s/QBm9fLTOEyKqQ2tE9TSJhxzkEDxjV4
3zJyHT2ZYdiIulPRx8JXtLgL8Nwk8s8tuR3ObL9IFKnm6OHvPXgZWZwvjUHaVGOCakd5exmJOuUE
2iZ887d6PmANMaqea7pZOYq+Z99IkJc5r5mXNdd0MDTd4fwpFXylJLYYvS1sBFZU/GSyvNC2eQuq
B7fCexfzCjup7dLj4H+RQVqglaJWGmu8iKORNhJLdQu/tL8P+JEG7uvDZGUay/8toXZhbLZmbFbk
G26nI7+Do+/6BFF1ZytXE3fVm7A3Js+bLpyjvGaoGpXWqKE23FNidiRxEsJmC2Q7xo0YHW7R/bI0
f9GggE7cxCGJwfsb4WLepMgf6A5qQhzTPIlulj0488UAohXPHubwiys7iPqrOoSiO8L3o6pJM++h
aJ1RMtrydKTPUH6yaDhaG4zy9DJGKy1NrmX8qNMTKyMq9nJD8JlR95MHtxAUpxnlGcBM++z/7/xs
iT9In/7Ye+qp4jgJ3sz4nornAt7csn0A7pwO/ogrtcG3cY+1pTb+FSz0Z7Ab2aYYNtLaLfOI3/hs
7CbnJE5SKDWvLpO6GCp+bf7xOijnbC+ip0i9yV7EMIICmvVHKwLWU4D/WKQgsxle85DGghNJzUKH
1XsRSwszTy3JDQVDh/9fErY4wyngNbCta2M8Z/E+71QWRNyLCHDrfykQY4m7AztUotFJgsm19E7a
r07qFrivkDYwq55MnYquZcbQ5PNHehS/zCsSkVupVXQE1johBxdjGV3xUEswAm7HyzsMhGKB85jj
XA+TcE2ezaaRnorM8WWvtMGqT9SlHUt8bHwfa85Pe/rti8FyS6Lc7PxIsdumoct/Wat/dk8CXCH8
OgnqyqJZ3D6dzq7rx4DGvA9Y9n+bJ8PSWDEfZaXCpdqziColM6ZtEeBxk6XM1CkyaNs/bnj5lY4r
1Cbnrc4SPW17spVPNJI3b3cxbW0jYMWUZRMN0NWNJq+HvKmZ/kwYGOZJmXKUazGytQuhzHLaZdce
lH7DA65iu4DXWpN9o2DJ8akZ5CRyZ5p/ohiu7yNt05eiNY07pPBm2o6FNcpx5Dg+8AKRlsm8ZWp2
b8kgfSYyah/W63QOQmQ0+cX119des+0J0vOoKba5Azc5nsvPKqrgrbsLyRQyiJhjE8yJAbJvCneh
j2Qc+dNZyCRpkO4JjCsCwsix4qzICVeo6F2mo5EuXaoi3SphGTVokksbuKjdV6tyr/RDFHHlOqzD
wjz5nPAx8KOxUxxfm/JvXnWeSgw3eFDsbTP1mrqGQvoyYD9PvkqMwihGFMCauwflqsQI9NCm2FyM
GvHtp0YPWC9HpH+t5SIq7SESm5Q71OPtHC5h7kpHfsuHp5dPNLJEA40OQC1UC0zGCUzojzmVUta4
ujmBSl4tYzHXcapukjR2iKUnfRvsEUf7RQInVcyOp4y3+AIwpdag/XWBsfz1ixxifvNuSI6aBSQL
U/C/S3We1xyndwRk19YDnkHglAjo277J7dJL6yLGVOe9PrEL+mOO5d5Xjp0JhjivY1OzWNSTuA+1
QTURAJxXXOSRLzIXfYXn+F1PR2ASgJjWOXL0nIkPRMLq6Y90SqUPYdUjYIkKRpqZAUGfnPcy/Ads
wOG0/HhmKSi5+GY6H6KQatGQ7Mm8ttgaL1Rjj9BbuSF2HZ5xKKJwhKZyxKbOQbDSFwr+a6UQ4L/W
EWFbfIT4AwENh/H4SSQIWFUe801/H+iTgUmrWR8sTM3+9yAqWphUwEG3gc923p5zF/MoM3YczszF
X4QMi02kNtMT6hsZcQ4gm97Y3pIgjiT8zEnvwhJt8RWDhQe+gOv2bGZ+UZ6A5eEnae83jqId9jMx
n4XrVcTx5hcp+zV7t+joAyRoiI/zq9U8nXd7IVH5zoA+sHmhMWRy5Pt7ZnqZKvDTRbkerRmGAL+y
FA3j7x0tyJHX2sPPSNpL9GaJJEkXNqCd4DcgHd2+CoxfN9OtnYWWbYLs1fFhvjG7dKjJ/VjY6jkB
cgMACJReFZDONciQiUVrLxK0WZwsehCngmykHNKHAYBFP644oUvb73mVGoA2OYP9C1Xq49G1aklC
78V7ZqIhmKzdkAszVEQOavSKpoBVKPWXU8Ml6tQPly5l65NntmuQSggnIfL7WIcyDKIFGkl2mWkQ
LQZJ2arOutW0mbk4FfSlUPPpOY0QdjvYzgZyQlMivfciNw22oqZAO9a24NZ5rCtd/HNDuE71Xz2r
z7t343WTtcfiSfgjRDqJ1enWRfH6z3QRdCqPKh0jg95VJtO3akM8nLn+6WZrX/XwABhW0n41zSW1
ZFRNolY2t6NFGMkawf9Clj0kHDqPLpEkT0e4HX/vAo7RgvLflt3qdjDQFWxQ5OX4OE/+VI+UdC2B
mG9BCITeSwV93t0aXN5fa5X90UBoR9cMoMaO/ZZdCz3h2kj6mBTToZZdCa4E1yN7bkwsBZgIfhRo
qzTVGGY1X/FrawqU47RfkGEsHGF+vbLmFzMtzqCCGgCvzPzg56AQvVUBko4+40wzhHcz0wIOSK+X
laYJ3/0VMDVd893VC4Ls6HBZIZFWjKM7q2ewoTGDY7JkHr8sEwvUVRx2GQ88kpb4TNPBT4OVsDpl
d+H7iYgMWSo2DVrw+CuiQJg1yZw4OVoTWvee2+Tywk6pRK7lKi/3W8ssDCG+FOiUoPXLyP9Iendq
RNI0TC/F/A1A89o/TrCircSg4lrPpZLQhcf6qFwplBHcQEpHK/fNXa4s5zocOt3DaKY+ily6EtpX
C1bYc4gtnRXl8+NDiztfIooVohYgEcqqhsYq/JPvRbdlIlXViQ7rNjOeOkTFx3Ties6x9pD1a991
PImeWyzwZgSAPc2IIyKDvBtCdnFd3pk+vyck5IlxAhQWktyB9Lh4yWjeAP8pdAJX2e1NOMPIaL8p
M5ZKtmH9IlbPJgx3iun/clJa5CZ3uB+SxmQR+sKqsssC+vPpXsYhR+vgBmxW/U/o0xWxckcRm4c+
WtJE95pcrfpPS9lapqvTH+HaHWHxzmxRPAkALZwapFiWyDoDaoTM2ZkzOXz0dULVZ1sXs/SoL/yO
WV9Ct+PFSYGXlFCZCENy8inxdieMK3RbhtTkzinQcXFXbFH3tdO4D/ZszlzqrKWZx6cA7GL6wSjN
WvnKMl+IjN7QCdW750O0pa7hzUoB2+nBajTVFgiE+3L6ITbfPXmOl85LmyqKH6cp4FsoM9hpKzal
de4zKUl5wsMtGzyXAY1OL4pzMHgsvJoeincyCscfU169PQ8XlE8ZlavmihE0tCY1O4qws+deViRi
iTBDFUisdGuO1NcUD5yfLnadvPt405VKwUzh8qu4cjX09CaH8mhALcx+RjXsmoLQ2XF/CSb8jog5
RQ81WPLt7ZXUbzq3kGRp07MC4PEJw5OhyThV1IcJXRZtrojR2iCXJaWYGXVXcOT5vtjgduIcG/Ck
x73syglVC318RpFzwBfK9r+reMTl7DlYBhBWuWtnqplGaGwUimjTfyLY2KKWrrWD9OHyzAWwwPA3
XTsCY45YtD8IWW6Ui3k9d2PHKSZZQPqQrnBQs3mEU0pxgh2krbz0Dlde6jtZ7GNw0RWLp5tD3AOz
y4Eq0RbYxtQB0PqwjmSgM38zqeqcGll9KNS7P9c+3ciUeROAEs06OEADfwrg7N14iCC8u3vyvDUo
LVo8tOE+d1DPP7rVMfMehjQvjce7uI7AuAt6yZbnGRb1VE6BvQ6SfJxPcb4VETNHYcadVhtP8mpc
8eA9IFbh0PJt9I3zIws+/lg19rbABwKO5uTXqjaI9TUUtl+R1hW8suis1PWCmkGnC4VK714pTkQP
Kt5EAijmRzPtV8SDL9wibpJh3V5b6KY6Rqs4cI0RjxV2jOzoyNCLjFd6AgUkA2i+rOOkurJgZtUf
B4VUqApRTdXbndsg10MqhnjKFBW8ze/bfkccpv5HebF+i4a8+GFxTdJJfDsrUrhXBlO9Yj7JqGGc
uj00/4GQQRyMq0zaBs0rjUsjwCsznao8C9OqSkWVQf0Yt48AzOABvMGEtbvoeZum6ZfMkL1nsfiX
cIA8r9qO3d2o54M1rix+QR33soWLnvtbINpo/iR2qkl+Z6mx5Ui+rDr56Olp0gPzT51lJSdYdYsw
Ap4SjPPx5SrcBP1sJ+eLOyCl7Zb7RuNEsgH262QvNiAfyA0Vwl6FnWXwP0VQuWHpVGrGEh6jk5Z9
gOlOhbSgt4oVtccQOCy+f/m6yOHXewqaslSIMTeKxEcFlmiAgAGEZaTbsLV8xWSkyQm5OefuOdd7
ImsFrGzaDVYAh2Rt/zvFEtrnkZU7r6b3AmDs7Fz7Aev/mxXWzNe62aPsnG7wrsqpBHwDQU1bkBhi
afTxzpCcKpz3e1x7T9C5+NbId6TgJKDDX8MvA5Ggb3idXP1mJb0yllXau5O7n8Cz2nkSWzXNjo2s
GHa++ce1ptM2kd+l3KPmyFg/KXtsqlWN4/DVtMLcI+6VItBj6WGDNid3yP5yoDdTAD6ftndIqaJu
eyBIAtzokG2ux6s7abfO55u+VSYt9exgmTGYLzdaMirhp3LjZWbwxjq2b30R0bp8bbbUqLo6t5fT
TH3SWqA6lI1086XRpuNe76yF/j9+gbe1DPdwBlpJaN4t7tUG/n23cDGKev3tAYgYiZVblVLlW7Re
C7aLHN+N5rjpIo8Sv/B+jETvptV/tDxPTA/F2kC2ZTVY4h5P+mZALrwyvwjGXRO7UWwCo0f1CnzJ
9T/baOsIaF8x8mWFj6sqSuerzt/2jZ+njoxhwi8xQy6BOKSWPjXFwXXyuWM01pN6X3cQA8wJTehT
vmmMpnn61aZadcS9OtXoOEhfXCmirjJazS5/2P9AyQPzrJ7tlZuNLEavIWorQjIy4aOiik76QO9q
xX5lzlkmJ/dqsvv53ZKYQ7MUFL9i966ebQDaQ9MPokR0ZoDrnDvMoizarrL9FznJ3iY4kuUCQnMA
ieegvjwbrb93estqN8WORosr+XUFtcyiQUy43Lecu7DgnA5AxvnWSPJfzTURlwRp3z9QBGwUeG/x
fDg9+LSBlvn87/nkSrKdIkaINFJkr+IUGUKixhsmXdFUphCTw7RguteWaaSkuaol7+iS4FqSkCfZ
JSyujevrnxhOav3y/XPoKOIu9HL0k6I2XtqbtfAkguJibdwrbeYBXhHiRHAbxRGGSzqPcypHeo8N
cTqRTM2Wmv48GntuIQYcfy+7VBHPupyC/Dd1xpZ0CIoVSI2YKFZ2rtbupGX8jbJi4FWye/QWApyK
Kl33UlVL7sN+m/o96hyQtG+C7EQtwQYOOoRCB7YlrRp7kCMWwAtroPh+H0dO/mXFRJRjvoNQN5y4
Nx4jNoqdJIYQKRVy/A3HrI8dTrSiqP1amFP9Kbzidb6klxoPJtM8qqlaq2bqLPtd4Rwn4EWaOXlz
fgKtC9DkXRJe1UkhjNkaNRKCaMAlFWUVplV2bILUdq/gDIcRWm5s7KyyyaNDIR/hILsm6H31lpkN
WDNFXpWlA9craobLJTDt692vWZFsTKUVWRqmmuXVQJ6Mgjoo2ktRtkFfUdi5YkvnJMMV90jxWOy9
E71oISoIJ3eYd9rvczxTLAY4RPJj1fwMQGphFWRCNFw0PQwRsEV4H3gZ6O02qtk1PJ3gDN8GpEvs
q6oIirFkyxFq4Cr1yILqkZ9r8uA3E+3zD8MV2I60woRqg3uCLnUQ0c6HcBSGPLC6tPI1xnDqS+fx
Nd5QTWfV6b90QW43hJSC6ElDN/M2QgrJi5JnnugVzGXaB7UenUcndBwgxE9/nCgF/uEWF2MP8Mcy
QwgN7zzHAm6H/pHLUtHQ1fMaDBb2xgeaJCP7sfJSTEBBXUBXFaLNDbp1qZ3aDMOiQ3v3N74Vevs9
bDUC1GvEBfL3lT3Z9RN0EMdMR9FSLWZrsYv3/Je2nz32qkOxv1rYeIPikIub59V1j9rcI7qBfFTT
PCySHNwB1VFnC0lDFXQIldRkZsVnv/0PIOYMtSleYjJgYACPtsvirxPB5f0awsgmaxKT9WJwdVlS
F7JAghY16+3OwB35MbhWtidUynFCp6razk1ondHMHnylgh9LT5vSUhu7pL4+O/btspKc/qNHxU4E
nVWqLmFuvZqqo7uWSeRVqH4fYmLuyVySaRcWNW/US0WaVz5ADfARPhB23Gq3ZcIEE5ovXPAwhQQm
FTLjrHNwGRJ2nM/LKbovbrZlHMiOtDbDgejkR144go5hZltKeGBUId0NUlYs15icwegVuccn5T93
P9a8IySLNChAFNLUv/cdsnh8DDoDFK+FyEEyIo+yOZkN4j793+zNf2nMHWx7jTyZgJviN5lOwI4j
8Nf/ijgb93rUfek6Etctn8XvqyZ33Er33wd0fC9QpAikxxKwa/oNwdHMlxZJxXcUXwLQQ2H0xF1X
XzUpQn8NM4z91yTxCR3OR/k+eJQ/z9ymPzrdNieK+4GIcKA26N6K1TARRAblbwbIhHRn0ryhGCBb
8qVtiM7114lvi2xX0htpsB3pOyyRMIdxuDBq1ooaeL8L3wN/w2GkOrTpcaHxjYhFwRG1tL9vQLJ/
X8uD4IY8wdP3tL1Nh6b05oYPwhrviO8wX+GiNM3KxgvxiqzST7MdUteEpYMXnz2fPhrcJvRxXS3q
wMmqrhHYaCZVTGI5vhaZLrZ+YW79Dv0kB4+Gr0OdWNt6uZoYTTG6iKduqxA3MXR6WKvmy0zhgWn1
Yw8IvhWyIUh6Q2J0iDPRhR2nveZ0lDrLa4pmwy7Q7CYPBuxu6/zqe2bM3QLRHAmVIV0js41OMKvF
fIYNHIntibNeQte2fffAfnLvQTQc83mgUJFEG9HYFo48Vd3c8Npq+uAQHtXHI2VJ6ZmUtM63HOsa
7cbyT38t35Fi5g24/u5/0OpDz7v0FALre89IpSh/s+Pm9ynEQT31m5BrDP3X2LbZaQCzWvcgnkvI
HLfKDcFOhYPkXXYwbAgaWSyBmgZk3vViqQ1ZFq2Jc2BAeL1el5tTeAsNx84iyhnWPupWsntT6TE4
kNJ6g7wu2IENkSD1egcf1qvLDc+eEtI/cN8wjhp4TamLwZb0gSylaljKYp5bJu0m+w9AT3cX6h1k
/kfzWaQeORF2P6R40dqAOWMpx56GlSo0HuzIXJSiTNK8l6pqsmKfg3WW01Jf89yczLyrzZeK+ytL
nl6zujfB8Zr/jltq3snbAIpZ1sWJM3tQhL/O+mXUJ1UR/qwaKWm5U70sIOxuGJSxcs8w89ESaYCk
m7CjjhqC+lPh3/vAXCXLfz/haR57JadeqXvVt8h/R0bdhhNwMU9LDlWOjjlcu41wsmoFyruWmJX2
ppRYYOqAFo8TFn2vRgZXTChp/hu4fhD64issHqVxZvBsOxXSsLpdil/ILzmBygi4IlwE9BdJ51UV
bIwXo2x2SOfQXICm2syqDYN4CjToEDbWsH9NiULcndkKVah6SHYYPixlN2M2skWmpftbnDBS2KO6
w+cFlglDDXcVVQhkwkerKkpeQbSHi5XEBsv4WX5wgmO9soHBQor6bw+psDyZeOgCSVljJkS/XWsb
wgD9e37U9FXfSJo1SgK6jXj9K27PYOZJde0C31egW03Ifxvwpw9Q6qCoLsPtSI5VR67RZIDtny4o
5thltXEXXXAqVBq4bDUs3K4ZTmmgVmlMnoxAscbkSNJ1FlDkHljsyX7gNzZ22cILl1ZUHzlW940N
m5uWHrKJlYjpC7DZ7S0fCEndQFTN7lBCkbgKj31aG2VmnHMu0Kp18M2vIVN8dE9fjaBikyjgRVlD
N0WOmrORYvUXojuh0ruMB1dt66e8zIcCFmO0ev5OqleWJ5e7bwARUy7MThyKuCCQgAc6xOZbuB22
yNx5Fp/LS+9Val/BidO9Wyh3TaO+3vLGsSGyV33eKwSCwBB+nYtYYsj3uVNeGYWmX4A5lk0gqfYW
wkkhmCMueou9jfz6NxmjQApR2XFJLdLXH/bHg3n8OB6U7YdxpWuNDRG9HMHhU3ps4Q55lmFu3u5q
1mvD0z8ztkG3YmkmBR4oEl7ZGJb87x4QIfWnU2h+oNJo4YZ7cZvJuyODuJQji1Z0b2NF8TVqRo0G
4qiOt1HGLpkFnO0GS0JDjGMYDLqwY7JUV+jHQBYJWH8CslEw+gr8N+5jMvkdJHRS/EQxcf4U/LCj
5d6ERRFbTpKXCWUyy8y0hRFuoXZiYI8Y2yOHvoLbataiP51+PJVuWTD+EAvjqAV4edAW6g60n6k5
bYovC+L5TNQyb5F1mMdaBTeKmk0jwwIA+5MIjg/MRSljQyYtOpHLarHC1T1K7W5wdFqyV7Flporx
otXf5ZPVSdvmvqiKZzZz+65hT0W/GeTDnEs0Q5O7wr6JIndcvegoBdK6gla/YGMPXv94GOQfYCyg
wy5UnlrjVTGF/r+5T/9POq7Qbpdzjuh1rOVmCHsNJ9VR2M+pBBDrYDy3MMxHmZ2C9Uj3Z4fvP3zl
T/3cc2XXHakP3QqBr0CiWpnR7SbxXupzUXOCqfcraAm6GrNLsLP+vYESWI1vMFniY+UleFRAkyQ9
Dq5yOB/YxTiZPq081AyZOuKwYatLMfvNnNTwUTqRX/VW2MA2+SOd1i8BqEmVQTNtPdxbWbYQhlvW
p8PDroF5X+OaWnlLpmS4D1USGAsxgwudSUKSrPTjkxupqqauzpK5Nj2qCE8BA/pI+Fslkp/FXW/q
hzYfjLchxXDW76pmZdJxl6Y044+98vg2RAImo+wv/kZwi3DgjeTceX6nsMFBXwaO1tkFabAm8DKc
jH9wr6qlxNN5VmLiOYhi6QhmU6lbgk3GFVAhtRWVT2lFnqwpxpVg9+H0L4lC2eCFiUpWnW7a1b75
omOm0bK5Wd5/vAARy/EyzZ2I9cp826OKxb9Qtu33N96VHQldwcDE3BqlkIMfeTE4dU8fLiEVOt/l
EKImDEuaIrZh/nxUhjZxmRglVgYoGHVG/OJBDEXAbHUbGH7Kp+5Rgjz96dZYDzURdkURH8g6JcfN
ZyQhH1/LMMX40z+OysqwKAlIDoUyTM2/qOoCQ924ORWgAT7771wpBUcvLLMGZEFbCY5TWnvA2HLL
ScUSKHwlom9cSladgpeR95DlHW8O/Jl49tjYS5Qf4o3XohJNkpisQKabQSYAJWNyZeG+ABx0CO3E
eswFjAcbas7BWAtvU8bMoSdn/FPzCZKXY5IUp42sH5QCSv0UJHfUtV3vW01haWsQg8U9TC+E9Irv
RLLZ5p9jdw4/4fl80FNqGbwPnlgk8PFPv+sZ229x/SUl7JFyDz7Um8NbZUFTWsbqqFS7A7cTauu2
M0qIbI3T0bNhtlLBcTpADVMFRq3++iF1lMuUBM5/JEEZH8t5U1Lj/QhSOdBDztd+KliGz3ZG9tT5
+5RLzep36nb2XEEMhvOgO3rnSYFR6zB9o6ohRVKnOeIn5sCDsEiewse9bDB9sNxB3uVMMVhKZbNu
1MXQcElRIe/bCPTDUEaAyXQitRf07jNgEBFzRyhqcF+aZ78ik2uXg/WUwIU9AhppQD12aPYeqw0u
KPYJd3Pkzkr9dF9WqkSLzLJ475oBRFini2wbw2O+JMZtgaHv+3/0sLhQF5sY/dbg3DwqVm3LNbf9
Wiu7e3wLUgbucPlKzHaJUxvETXpjO4+Ujm3RXzKn05K8lD0gAh2UTq0y3D9TlIMdVRfbKL3id2rl
8KVrqy8OuRXvVVDqvRr+LVoMeNDP2t5PISIRzWGsnDHJ4Vrz6XSx44NNivG1Vex21ASK6FhJuZzX
P1tvfwvpEbmu0wJeB5NJ/dKwI31m7QozjcbLEOnyNnFelc4u5BUO6knbqLOMjdI+AP4WAYFhVVOG
x/Tfb96mDzO2vnurMFmjTLNwHSWAp9djUKTKUPXUpGSepnIrm3U5T0IP/rlBVkc8a/+B98s/CIC6
A9OlRyGNCHdu86qE7bbAkdUhJJS9ZDV3VPnSipO7oY9Wa7zUAGzVX97X/4V4O9x7VsbV74lVYeu2
C0Hu29zSW49L0IgkLokAX26uhRUJ3nDlfCTHLAZ0d4oIx8WRy4Dz1pHOQEtY/3O8wwN/rjP8eAfU
yJt1AEACM2PwJ5EueSqOTM7UR8NzWERkcUQKLqvfxz5ffC96DgsU/BPe/S6usVANwaBQB4e8/wl0
09Zij1zUG3jy0/2iI0lu/BpQlF+TAmfRFESjAO9djcAjnrqWyf1a+YAlBzBM90aYuIWNnyMwGaI6
ICw8nqg6UI0WN/W6ioiGWMK+74bdK6bVXIo6yoa8dgfIdckaJc0Mhbr3ziZafUN1fCQE6YNDQdQC
xPGhwDdXpPgHbm0LW49xZT1j3mzwxSoSCkQj0EcmPMukr1/+XY+Sa7HQGZwWuR1UI6H48YqPaPXq
FOqwod5OtVO3sFHVApW/DTW4rZHyGqFyqiTVrDV5RJ1qSCASDHudU4VtKUx8irzy2P0+GN15KpKe
zRKkrtj5WKppx97Ztu69Hxk881F0GhKraVuZ+/BRGurTkuPOfR0u6xCgzbJuMadTarurGDczT25D
umTGhHe6YZ5AoVIU8udNvUsNcRC6if/sKw8RPOExzpc1ZpwkggbJiVv8qvVaGPFLtYGMN5zaPkvD
+wSpnDbnoV1e4PUxrDX7qdml5zkO0ZNioDAIhv92zST/xy17gdqNn0LKF1U34YbCro/QOVHqYgF1
O9SZjyFXmlsrqwrQWRO2mX8TPAFcwYDJNSKSgCVcs2dUWZlQkFyoaLK4ybSQqI6rLCmjp8l8Bcbx
jSmG1DF3JpS/QgnBGaQycq5AIFwZVTuQ27pWa4F9SAtvdwI31pPZZEsftXUbx/szHpPwqxNKoxOt
L/n5N7vXBrU+g81mhoxyn/DC5OyMkF07f4Wn0TWpT3V3w4mIXesVj180MDZcFbcfXOL1Y9/9V37H
gxdVwlZFck8+99OSgqnlo50oR+/7kmIjzWLcS3paisg2goys+coCY922MJlLuFGm70Ohn5ivCGol
xP7j9XxrgBugzllNd4MMcECAe95HDItC96z2kxiZFlXCsCN7Dr0m1g9i1TVpky0aRG1bsFGKCimP
sdtk87INPKbr3LeVYEhCyT6AZABlZKpAe7wS3UCKPw3WvIx6zJrzQ3wXY8kSAYcyu3GF4JEXoa3Q
NnNXkMrjReaye2CicXeFFmV70GDVdMYxBt2VSadERB7OxEz0969RCcwrdFdXooIPyYGXYYoHhmt/
FlKmsyziVT6/husBZbCea0+SOVRIZPIbtn/adO+nKkLJz8s5SdyVYeq63RaF5frwGvcUz27M6fcJ
4kD6MydSMd5M6bJadypHm7mqmvI5laO8/KpECcLQpETU1uGk46CT/yk/kra/PgtLXtfKsymAEBlI
UxDNpLgMZq7GpIxqQTkLYASEj8KPvK6t6Ss8EHtAwjnO4o84ue7HdwlUwgrWcDQYkqYSh4UyTwon
Uvt7m5JfiZodTry1qVPtp+n9NRmKUVpEJQW9GOVqEzubHcsPLc2cmpxW7hsEabQwpVihkAcjvG2g
i//K0AATaKbuV/fm3SRUzW81k/yOM0NT+1SFCsvyS6q1dSBlLXjDOSbagHOynctOC16+yebgkpit
sTzHuT5BN/D7cP/uM8UHdOagDP8FwiB4TzgGSAX102XFk71X4Dr20yS/e3uKB6/kH49Ng2uWzqlx
4J9acS5JJTlgYqicNDFSJI100DSPCHoWGa3KGxczur2vYIFe2FIA6VFtNI6BVy059V+Dh8kPbCL7
/03h60MJYVahkuNLdefrF0+/DBAu90vvrfyBFG2YwjsiDLOhF8+faelJXAADfpx3rynqU/fjggw5
4QElAvq5NRBAQ3F3L8p13DwD6tZ0gieUZ6fsRyFXQQXR+y4qbcDH3qP+annNU7rWtA3oSXL1p8N8
AJnhLaVsXvsawz+EfLO+SuVQ1BaY7zHa6ogSKiSW5Gkg4DgVJbcRCQACest+uNUB/HTt7UPQx+B1
90Kaeg9NNCB8Pbh8mc7pa9IKvm7mhNP8aDK+zC1tYZWyjBl18JpfLbvSHBmms5+3Eq+UHjYvC9oi
UPuO1K9r2ANISHreBR5shhNfYdolly82q+w4kzLYlfU+B37FcpxyLZ/BF0qFMcp9m8GIuplENqLe
QAkUZD4PlkDB+4pm9pB9A2euAUnumbh2pBhm91JgpNkdC09tGoT3ahNzBK4MPj6cUZH8nKxOx+fR
/YbXAM85bIswGRNQ7//+WX33/O1kkzGIaKms+38tvyE0/7mzFQyKv/D5hqvAd3pikKp/CDwdTlSn
6B0AUTeh3UVqVd7u8Quu3+e6cl+dX7q/E8ylAKDKzqqEenH7JaG5cHG65DndnwW4LBvdId/AA3zD
XhXJYAAYNX/tdx2VcmE3AilXGPsw2ZFHXP1aYoBxkA+xespp1HgTiWwklTV3Dh28mP20TrC8rV/F
5k8GroNJhKDf5xZFeU62O86aJYsbeV3ACtZYowfTUAi3UBtIkBhdw2YfrT8yVAmGIUgGR4tJyjdh
LBGkpVfJUHqs3Irl6jTxOl9p1W1KqboDcSbgdN3QDOu8g0WPu0aoiS0RV4pu08YABflMG80IQhMR
Auw2YHcH15TKft+DsbnAYxI0UJAC9Fx1na4ihikvupx5viLpJYK3s1kGWg+PHQ3xyyy2vnrp0QuD
3TAYtW+HO66a/XV+ry5P0XCF+G14lbquzmt6iPcllJiDHG/nf3bF+1l2ZSC4jNxkHHCOMxmBuua5
Sm4qnZNeANeaK/jrDv/ME/Gm0VOfeVNG0XRaVLtbMY5UHOkWOmmRxoTKNSN9U/Fpd3LGqCRKgoWh
1z24hJrYtg0joHLH4Q69lB7rtmq/Szjw+TC1Pv4PTWlvAzDB3hQlR2B6VAZAh30oZhJ83ZsAyFsw
/H5e7mFYGRurUPmE/vyfW/Li+FJ6iuPt/NEwg3o1yb+avD9WKyGjgtLiacmk4vEcoCOd7xJHsASr
Lq7OSZrgtHiU9nrOu7lWFHkxAAQURQwbXO04xaXn535oQ/FG7fa1jhv0SXGRnIkg4kZZmejir09P
274qPu0wFx5tlwYRCo/KrhKvBfkGEV7kuCGClUx/pyDISK6wj2jS/KhpEL75YbdwOnLMMM+LrT6P
MHU+PDphn7kB5B/J11lA0mNy+pQ41bwqXmVuihg8UFHGI8X6EuPSaHMIwuBsZozli9IGnfcCKM6W
vh114T01E5fkgFsm5XCpMyf4Ua2y+d2e6QcuSvN6gmgqYA/yQJ8M7e4zgDO2eEbYcIP7wHagHuJj
rHVrf+ARPOqucvOMNQnhZhDgDo4IWIgnurm0K6YaNt640ywJXrmswsI4SnEgZtyQ+ApchkSSFbcD
U5uOdWYVVj/IaKrKGxUs0YpsBlBnH18QyfOxiv1Xn7Gyu8kIc2ecSG1KhNQhipP95bDs9fWTfUqM
031OssO+TLApwIJy25yQigQfQx/qnl4uGMjV8PschR2iVi9VT5wV++ilt5US4ohd5MsRIBn2j7wB
SrI+upKSWjCYQV+GNJYUEIizF8sSOnzIr963QexyPJrnPBYaxoO9jyN6xy7rEZgcGFIVHLfXQYu5
4goxKSUmFbYKUVM8HlA+KVm7nyrk9D+kmwGTCpyc7/63mD/jhfDFwtiuuWLDib1aOwta+8qjgA5O
b11mVKUPU+kZ4T4JJUOEJwoR2RWBPQW2nscIThffEF8JbrBaPAfQtzCh36vcFN8yXmbDAAKw19Jt
RXzmS21VnpnYPBc5lNXp6O6KdMF8Z9Ey3Ot4BF6lrijUdUYDLd0QszBw8FhPvO2DkgHMI4jMtD/e
Z5fXruwNoTMqs7OuP+kOIVlhkFJp28hxv4wj/OjyCsMKRIO5m2x5eAdjM64L+8cfoScL5LmCZCFt
BR1+dzTQizg+JqLtjuYu3a5J65iHV60VkYMkfc4GBUVHYzMc90QGUNWSf/2mK7HPuoPayJ0WtmIz
47mR0ogQj94as08Ed1oh0JDe20XGSfvLHqogvzxoj3ZPAiO4Fsri2OS6lMeiWC9obvxi2OcwBZub
0WRQQCpMFwJOzJvkPyaVl2+dPFK8TsApZmbiQD69okKZClBq/x6zDjTBV9+7SGvtKV/pS1+Mv97n
8Syq4cIlxzjgQlaq0Mf6rnjh7XOO//HiBcHt06RnAczc9XgG3bmSnMVZwMgGbLfuZmybt8qt0jTH
0clHvk1LdILJizMjR2w8XtC1uxWL6nmYAuW/BeW4Kwqy5bz2RI8MrXJlVb3j39PO4KT1AmNzoI/q
9F89oyvs5l7Whj/H21RCMGZLwPh0ui1XWltvjJfql6g43P0dzb7KR0YUFvUNYkzh0E6JcJoK9QHz
9KtEx6ed/sLaLV7RUSCAyQlfTY5TEESIo86r5miAzNHaGLb6AzOfqVCUsCHLn4O16CKEzd0HxU4I
J+U0bEf7GbHpXCB159UBMt3KlyEPLuHaQMhdEcXfQMVURp6YQD3Hf9h+RKY8ye6aUvlrUQhGCW/8
CYeZL1uIvty4Pguz5MO/e5UkPUXAm+cX0q05+Jo7EKVNj26zzoiHOsS0p0qwmHgfTB7XPHSLm56Q
2Kheaq2HGLWclzeVsIlkCnZNYaIj4kSh2Qv0HI8IZscNhNNClKEhhnzMhwAguiqplxBk3skf6GfH
DeNa1MNYmPh2JZGYZ/sxNrMGfhVJpOWGWIY3oVj3PE/eG76m7Jow7khybBoAulToCX+SNSFrXoV5
3OxevP/RIDsI6h+4nDgeLbs5w5Cipdqyf4vsglbXO8h1a0/fOQWjou5kmWtb8bSckJN5Ql193jn2
bS7ThQVsQYPh4V8x2YiA1BDtQuitoeopIws+f2ZAn5PkG2jevytpjJDLaZgzGPB/F5uuTzSqhgjc
xTlWJyNJJc8376d821SpIMMvF6cx5WjRCZuwtWLMKAJ8smFLxziqN+zS3B+nu4TKb6Ln1I1Qikmd
MRdDpNku1cC9TtrrC+Vr2nGgbBrbDYpW3lXV1luMB2KfD0Fw190VQ8SmICqqcG9j8ZyI3qHCG35z
mv7y5f6n7gmMik+3aI3Tvs34RpyMmAm9VVLVp/rlrnDXruYnOMDoOjTMrXhGDdoyQU3RMByVTCiN
34ycZXSREsgpX7Glao4PkfbI81OuZ1ZgQw4IC0pWTPYQqkYwZz53vcR3SR/ZXHv87XnIz6aIuuZj
OUHs0MjORuYwxN7ecboVBfSyGLoX8dCVEdhI/1GBYn5X78BrPszH3dwOHIRYfFVmtJ+9UakMHw9Y
SODx2pDzNQIKbiYwer/LCcS8Uq5EtyoOCVqiFo7L5NEhl9kN2fQX7Dga94f9KxR1ObR+5Ukf91XZ
SygdHofwXbcEMNdTNDO43/ViwuB32LMsbdNgTAXOERv6l9SqU0z7NEt/EkhWHka8e7XNJCo56lbM
9ySL+0UCUsvjdYZk7exdalbBk4vE0A5AOsBhiqutllAjU83gW85+GbTgxI9pDQtr3JdkJi1vk0dU
znc6SQkZfXlZ08kakZTkRspzxbOdbNRB5820ZeB1k8zC71EO2Hbqjb2DuvVBU/eFLN2FtyirBh5s
l5tAAyRRsF3Xxiy9z6oFRpH1Uru7ko7OEKD/2aoWFkkZ3y57tUGyOPY10rEorWhl9Q6ENzWcyPde
UG+0mZ3jHa7VUPd1AXmCyjp/CZESBXNSNFth6vlMKYVO+xxt7XyDrpBWqfazQQNHEi2P8ynMrAmb
rokzeEKMmYQB5eMKro7lVfABd3/GfhO1i/G0DxhadqkV7XkmXAH29hGe3T0GG9ROSgM7sxB1W9lm
73/n7OOHS++hNT/KvezIPuSc70vgRdX7WI9sosf9zzcrBlMcNKDtHsltVekKCluTsMENfNQroc9c
wNTDKIiDY4n6vg9FSUibv39e4hdBuJwUSPW9ElV6ST0rw5I0xDX3fjygA2f91NwLFYyWmqp8jZlS
jYV8ZpMoko2MBP5kkA4RWyfQjtgOhBcZT7uRLe/Luit/105aFzNEn71q7fckl9QDyIiQjwx1bcX+
aPqAisOf22UYVJss2/btKqbr/Vjp+mGsYiGNQ3+d6OfN0/q8v3gBsEbX+EmGjkUPBLFUUzCQNZWQ
r9OIS2U5FyWdS2fA+4Mm/z7zc3oZXNEglpPRiYusfUqs+1ZGBupSdvbYf0rdYj/jx2Mvkq0hFf3/
xQ1HQUFfxcIopXH2EiGLTSvd98Prhayu2em/v8mxm7Vm+bPh/8q/BBscqThv/t14+LrocpwlkTsl
XzztINRz56etsH2aW3FNaDSB0sogZFOYp7jVD5DFCNtZOc3kJPY+I+OMwXGYrn1SE9jN/F0PNzgY
fvbGEt1jX1+reLnBPl/ehXxtZsyOt9LljQTV/eLlzrz0KHVKjmAqdQI7s3uSNanDJjPg/BqKPL2h
LqC1iQ0lstr8AarcFXGuMRkqOIrUlfL/XB7IjQ7AyJtu7iU/j+7mu3PACcZmwDzBpKRCn8kYEXH+
VZK3P8LHCiAAu681LAl2zsKtBvzM7tzHBBfZ97JnpJVpjr5prT9yaKKmj6GeTH/3QYatslgXP1FS
THGDyFb8lOpdEicOiW9JXR/EmC+kLf3+z7JNh7NW9pVNuixgecSPXduwZgN8LLUbGFuAzVM/2s+Q
rkV4d+j9rRyiAdlAf2X4MNgG9n9cYl2sidoEwVpS/9j3WwsRE6wMVqJdYz+gQWx1Cn5gC/KG1OCS
pgxWfjQuGtkAPc/YymcPD0BiKCr/sGmhgQjEI66ds+5obo9HjBwCIEzdCHpCIAUKEoM7IFOZVAFP
N2xSRLFr1YOF2xfcFi+UUbEFoRPyN/iHd4CIuUmvOiMgCy7MQYVBWGm1d7Ffxj9sCWMMgCv5hjCb
JsxiS1gHm+G7CBl6fGNuG7eAPdmE/uw0gxRZ4goF8ELMlkk8Ihao4qwwqc+U5jil6doUcJDV2Dey
IynqixlHIRTp/OFNcKJzInJDYuGDBqT3jbMoYiS1EY/o9XZL0MrQUXVmN8Pwaf3Ua4UwXO+sND/w
DwsBQsi8EGo1HF12tJNrKBN3jTUIFZmLiLuHPWHhZea+JnZE/caLNmbmZ6u40PclxR8/v/5cyglD
OHtLPyPv0G+Vphf2LxbzVTw287VgAzVsU0Oe9sYHGirzXShYHe/7xTH7MvK5KWPueTS0XPUA20s5
io0IQ/LZUb21tvbOGC2LMLBSTUC0sJemlFqDsHe+EQzLJqb6LH1njRPLT0TNBpYdqM0a3NPfS93F
+o/oPszCORB4M3inC7SqVYvhO36Plxp1zdR+clrXDau50oPBDXg8Rrt9Tau5U/AJE3qCwXV1dMFv
W0bu28oylgbDPJuSRJnIeyh4o62MgqKcUTYjtjUy4CDj1xgGeH9taYIisJbfq3EFYehP2q+xexr9
dL/ENrgwOPrX5P9EgbI6+UFxyRnUYbiN1eMaiBDXnO8UftbIG2CDE+JJNo+JDKkxD2v8zkdutnaO
HcVpaz5JRR6zxPoxigaByKVMts1wwMZY4GgBWuUQo7W4hLqw92GG9k2v4vGz2kF3XywdhCG+4Lm1
wzCOXuj9QhGCDvE+Z5DVYDBfNSs2pi0oPnlL/tdH4E40hfm8oz/DauxPnuomT1wiZJVBGW88qVkg
PldqXc3A72yrtHXxDFLVUXiQUUnVAcZMiX+82f1RH0GZG4dcelEsDOq/2+iSEa/blVqqHPELJx0x
2BXM/4WTiXBiehsZvMh411uMnaCE7bIiTGjfCDBNCXHqtPcQBh+RzoHdPfz6sScUUIQ3rCiJSE3y
c81AsljUl/eg5g7QbEEsEEsYtbeYsekQuXp1hsLRl8aMIIJP3KC4WQNvgvm6wySl8PeEX+FLXdEu
g4S2M7vN2K1lK4WyYVZrtgOULiF5q9T/u8WH58gj1tcN05fMtZAoP5viv+aITMLzW9dd1/Read0H
9vqbLlLfUKg6pLLocjWEsotVSRy6wwELu6K1mEQLA5otESLNt5weD8+pWsvqUMZCkknouf1+B+eA
/PTBTKZuSr7LyXbcjT5cvvTz0Bg1nlpo2tMCx6K/Psd7Y+QBExOdVvVKDRvbOl/3c3okaEzzBJ6T
UmnbrsWkUC68ESI50A3ZN6Z0J5w3j4MQP5akNdcv27zzDlWTqLgNrzWRg+UpS0rSLJufQWU0CdgX
w35BRoj0PMcOryL0pg+6/WLY5zXE8NNPmhWajI/raXGGOr1/mW7IuP6nk7q6u78mnPyYOSBBTk/H
HTrDrEM1vzqXQ+F4ZDfhapQHOmkdLVWrYY1hiGyW63EfqEMzo3i6CpHQc8H+i7ZPfHUMJQkA0KrV
MXKaS4Te+8IZc/tFMtpMEBQRPCfgdqFFmG9bGLRAVySung4MoAZGZZA2NaVIqK4K5TEXZnRVeISF
+Ph6Wh3788nOasYxoyeIbGN6jMHu6lvb/GRane+I+bZUfryuCIFhcfxfnTn9VCvBIHD73QvEMDSA
J9MmhewkIUvC5yhl+dwphHcWJ6VjH5bXe6PEf54SNYQ2DnFIGfgP0RcWcE0S1aq8eSO7SUTwSkqx
UBLbmhE0FTxdg+z/YLKjZ9spxdNrGh2pqaN2Sye4MQJWhQLyYs6sui+BnPUYxtUJEZqs6efdExHP
l1eBo5YhEEaZUIeNMz8iLxsNCBq6vnm61BTt7F1T8c9xEoArxFbxdFmrPnCABZCrq+HwAmPs5Fga
2SZNahQs4UrNC5HkvkoKPY3ayLPrOQ0wvFL5XTPnZ3EviaFkDp6UEJ5ucVuMff2jMtYZKZ0288c7
DtdEgZM6s7GMYHcGGbhBpgM0PE+RHCB3zqOnqpZNwgVXEswJUF8WQExJh1/ByUk2EsQQNywjXbOn
lYUIj+fubUQC1OwW/hQyLj3kFGQaw2Zb/PBjZkwjYVSaJ3oCTUNAKk7HpNnc0dvZ6zomB1yDvZdL
JO487VAzqQ/ZGcEcoLgtCAbWx/1qlRpEBdll7yD8Dt+ML6/Q/cWX75aRpUM5Uc3qt8R0w6pXkIdy
wqsWiIe/+gwNMKTt+njs75Z3waWPO52AfczMOaiNMJUcYWbffyrpf0NovhXA4nK048WoI9VXv6ox
dBQYlcfJkVwuTJfIl29LgHPXDIS/nFMd5auh2OC5sAcdzV7MgVltum38PCSCz9PO0Fot7sec+Bs9
CUKwLRMEvW5NiZBiEvBq8SBgQM40hR2+VCcUJo9GJH/yIslm0ALVNUYwG6y7bQ6FLSVt/YlYdhYB
EVFvH9STzYzjEwHxK2v1FqOXw/eVLzyMvNN+L+zWTSYXKMWAxgZXAqJL5sKp9yQlaIirJUhioagm
dYcsgNXfNKWSu7jRViSryy1Q8BAT7kQuNpnT6SyiWsvhbhDB0uKwgwAtB+bmxX0r3kqxMxBJWS4U
mmGUV80jZwZyxd9QwzkFH6COg5h0EbXaIM9m2VGoQhDKJGVGs7Hd5p7SgIz0+txNx/ODgH4GjHEP
icfZm2qtOcs1Nc9xmEjYaihunDszHH1ZjylGF4fGtzyrUu7Mwd1BOVPME6vIYEwRa8hn1zP/WZYu
pNq4WHpzzRdeYzcKw2i29QaE6472V7IdEoVcRImfBCO2kmaKeCkB9nmehOA+n/61CWnmbLpMrxUN
HyZr1SIr+JC27zCocIRVibCv5rhN/R+jSlJkd7o2P3kmdhYc3S8W+eOQ5AenY2lB1aQQpTVM40zW
OPrkx08dIcBDx977ZDlJcP7KVopABzvrfGcFBVyJdG51EVwUePMcYk/fleC8MQZ/aCPE+zr7Gdqz
aKFyFUIlvIBWgr2nzUfnIGZhiETaDTnIiYRR4kWAE8Fa7UBzqCNvEbbFABNklPVbmh8fFTSvDjeX
DvExPBiSvluFcJX+oG7ZFkSVdXtqc7WjZZ6V0KdRtRkJhZ0TrbaUDYRQEjwPzoF+ddvwzGzoPIjq
8FiFAGcV6hPgcxxTTmKfxIZ7LoNGwbQwKsrKznvXQfcEUt8BiiiVyQv7NrRbBAPxsu8a9TU1DOZ7
LeDi3EqJY+Cxb1R6KlVAGsBXM/GpoYy7XHxWIUrbpKdttRTpsbbB+Kvk9NPF9HUemVM8yn2cN7Bx
HAYrT2hssvXQTk34fPFdXdPxKospgnf40lOHPw2zU69ojwDGZ2+o/yFxNHvvEgCiSDkKV1ui7sCp
sVA4CnPPtEqkk1HMIEKAcBktKZgsu34VZkt28t8nRaGNrJiYxnUI9zzv2MJ8rhd4VYG34R45QZ9K
ITufwq2vB9iJ3tQ4C8zWHSQc3jyV0DXN18Ma0MtrJlt2s07Djc/54YDKhaLgbNWR0zYYvduV67zN
zvMy1IQV5BnVFZKwG7p1H6b/dogCpDcwGC+0XfU+c6xG9/b4LOJaN6K0Rw2AbaeVhu8CopwG2C7F
xj7YbiHMM23Ut3jyLb/mC6U+aIB8w+HHsePdHYx1eetLNyIZHMxAo1YV1D5xsmqPYaYxk1N885Gl
yeVJHFnoNVqNr2C94egEg2YJHVuQnyKjgOa8kElvSO+0m7fcPT/PPpwjuiTW6/YI5+jO6VaVkrTz
TjnL3cMrKcmjmVAnoDvR6LpcAQTQgCugTg2I+QkHDFLf3UR1KPkQaw9NfZVND3MP/dfyNfCX+oPw
3zWZEXT8bPFuPtVNoXgh7fk9fVNlq2g5aP1KQOuCKXybIvyx8eJhur8wXbFK3tOQ9pWDveDFrVcp
nv7SpY6JKoRqHtzJAHomCRDu4NY9WrhEkaWTeVsHEV+uqfxNTDhcmQf9OVd+6iFt+NJhk9FkmIhb
sj7ogMRVzC1v4FOqqj7tqOoeDuTC3vVYx4ezJbGIcAPO//Sh8Mz/H5a3G3VvaY+w9m8EAf8AkCCp
H/p63SMi6k1MXkqI5zSuiHpzFmB/EUNaOPCrwDF00UpzfsSQiclzwen8pOCxiCNQM95jtV4QWpju
YBJ+FkaAyXCOP+OdWVoa2d30YBMg4AypAUSCbBQbCamuOQIYMCN+zXUN+DPs8mMjVS9FwcBjb/ag
cD42YafJeQ3MiCAfOJV3jgXsP5a6tk9YUQrtTkt+9s8oQcCrILa/LcIAcH/V37OewicDfHEE0jgE
+/Vlh7x5Y1b5VqHqeQbWAC4nTc/QH68Cslq6tFXSRTDXEjnFEDBi2iT3QTn2/uoDHxxKKNoAdRlD
uREvG9bhvT4SGXmN15vLwDcXEelWei37+mr973MTGYqVYqfdTsXozLDIwr1Gj/r4jbUHFhnZDLpB
DEwI9XJUkfTai6YZPFFG/BzPYcOky8fBnjN1h/6fK6k6hJdYcAEzhDYgWfsoRk4j6rJ/g5pCpori
KPnC96d3eOSMAunggQBwYDpOAqDM+gsIZGTWBjd8ZtlYCpPjEbPFFD0ifACGIS/gRY2cWx0ttMbF
ialOZYXUPwGry4qbxlHpZbdjcqYfxHl84IfWdo6vZFFDxNP7u3CDl1HZrf0KVqXYpOgzSu8NT/ZI
qn8bK0hbGylRDJBnT+m4Ji+y0P5SlIh9j2v9wrrC8t2XfGA45aE1aC2yGJJhleLuvLjExa0Ao5uT
1XSiiDdf4Aq6ByJEIpoZZFKm9pxFUPt1IO/KajYIx5zRpbyZ2Xd4SXMWf64yg5ap/79uQ2D3K4e4
hmMW005BPwoVniHswN6Mz3pYKCEU1c2wmU0Y9iUrf47jJVcqjAO9OgBWV18s27kH1MxCUZyfvxg4
v2XshTa7tJh+0Sojjd3Oo9ICWOszEXSx3U06IFe8BldkGKwg/PYzGtsQMpFmkCYaFAKVkYvIv/G+
E0W/jJP/AutVPX++rIwEHlP8QSgJrRvojzoDG9yGS64PN+GmB4VVbdA3QUcAs4wD4gUX3qcYKB+W
fXsBit1HNOvUqjVoqZvgVOHq/IwZUfzpKJDjw3PW9mn/PISs3GmBVVlG39PPZ7piSmPXd8/Wwtfb
6iqyvq8Ar+pAPBe0yM3WbWvQ9a4MNUA/XYkaHqsVNxyoFqwZz9cjB1c7nrDku2Kcc0mp15qOFlwj
/Gm8d8yblGrzqTPiu4j1gzzkEHrXtibaCvoJtGXScYcnUQQ8lQMWkyvAxVb8HsaOW2BvB56DNZUA
t1qkFqOAInod8rrBAbOC4P+9cu/0KuYyY6gLCpqKcmk8DRzY8nx7Lc9zIbufUVVy2nPILPFpDQ6r
GyDqfny1GBlgq7uhuXXz63v4eiBTj/vYCsHP8TThc4cswLW+rm2xrMRmk6KA2iacjHVO5b9f97up
H/1Dk8TmWQnpzFw5bCYeydU5cpeVEf/mHLYNfMjji1/3q/5ha+ett3DVKNEyl+HAUQOJX3ejeQgh
/IMHZY0kvLqnInvh4Sir756JqxwmIw1+cGEhpbnmx3daB2T+TCO+vutWwLasDSSZ7z6CEnmUIKlF
L4KRquAvjdwW7HWv3f1ydd2pXjkEVvPakcRO+tc2CzfEiV0FnSOzEaQNXdLhnwTVrOo/FRaVXeL4
eBA9KmQKQFzsBLV8i9DblfcFPyA1MzCU1hdgpGo7azyGr5TgijkdJgbbFtr31ZIi5swtJXKc+1c5
ACJApe10s5qLPaKE4h32cyIHGZjvkmysITHTAHy3owRgVeeaJdNDTeVMzFw3H34lBKpC8vADD7vB
T3gVZsvHgXg21eSOaWX4qi5GkznTJkIZmq5ahIdQy2VLBSaPLcdnK8YHNysg+SO/ufB0JR0Z68Vb
T1sKIkmCtqFL4D5uXpzrFYXc0qZY1RYcFIYYhFsc7kqXkdEkYIvl0LVRJxnS4BBxlrDgopP94k6B
q6G8Fl5sER0g3gxstJVt1yusKuezP+ZAYG7ItJrP05lZlO4jFpKcTmF18RcXxbgyfhcuNJ8wFwiB
vECqzY6IyZMn2nFbhsYhybWvIhVYGYqjXa2sKcPiLX9EL7wVWEZy4wES63QsVI6M3IRIxZyayX6c
xef22Edhr5QX8toc3UOiN29CMaBT6lHGqnhZYmU0OQpVu4KdqtV25+3s3ymAncc0HuyENsL06OPl
LntVXA5KVHqD9UR+tUn8tQmu5grS3hQsdCl0Bhwc3DmGuJjUC+k7y8ADY7HOGbIa5LipxhbLYtdh
us4LsXvaD7EItx2ouF1/gWs/2ihgI6NH0zOvGv0bYz/aAe1OZIapIR36eUmnxW4Qskm+LqhbuQFD
t0SVxv3FxLSR94SysO+vbSU00jxy0nvikzX07Fnljew05/kNeVFCIj7+uQs4MIvhla/ivS43E2e4
jhDfAl/XLs+HVB1e60i8cXjhSDTKiklkhw133HHH07xk0bcySmAJHHp49mnJl2b9TNIARo7XPpDE
ELgAR5DYnir41nnV1ZtCVfVQWTA46firgGifjnTGSsfFxmmvUsVuiCG73pS2uBlI/Oybvj6z+Jlz
N6E6stIbgGzeK0DNdku8F6EW42Ulzuyd4swVm01iqej7H3sQgt55ImiK9YBdgU2pHwoyr/fYjV6Q
0x9nMNh02E/RHi+WzAVxjH5beR1hGxHKEcGou7I2rL9pLO6LS9lgOZ23OFnjdX9eItsehlsj93ok
RHWza45F0L0XpNEZympBQr2Yu9S3VKD1cfGGoOMon0nsb+f5B2Hy/sWAU3Q26WJGtH/ec2DARi92
zBp5hHcZ4JRZK8FxI+xyc71R2aVJ5+EICRGqeFXSOGwjRofHN+SC7A3shNtrsDMoBeRUDcELr6HW
wV45+bGNCGggFKryvb7Jsj4Pk0/k9TBH6nJuy4Y3whtSgaVUakQfiRpCpezUrWSbX11b97FKOBqr
VAwCxI8Ijyp8tymeq1SyTcmk/RaIu3hrrhiDcVLzHEti1yn5RteYlTOxHZfJTx4igvathmjJF8W1
ejTIiQBgUjUFd8VtTtCa1y6+0Ss0lWm7wBMYuOzVCVem2HTX6zZIs3zs0pt8yeTDFUmwPNYc7r5Z
HFYTdbDw5RfcY/eQJGL+rU1FhSoD5Xy3r32WSFzgO0LVlBrVgHZ3I+9VAFLjjrEViRO7kWInhcGg
OnmiMYiElAOHfTiui0UmlU/DQvIPkDjqJaPw0cuYUjBK0x7E4s7GD2j7B4q9UbEjM9pdvsPAE7gr
YOZjh1Dz+qBN2bFsb6Lh6+WpAlzr7rjhev9617SZE7eLLzwpu6jNHN4fX4Pc/39W8PJl4+b5SgpX
MKf6w1GKrYvrTKTWuKhCa8CpkQd9Hpqw2JBifKmsy3rOQBDJs1oSpLnD27V+AwBaDVHBSejpap0E
61VZMr79USWDAz9cr+II/zjkQme1gFxtZ1GmxAaNmeIezEDZYIDZR74znRjDGEOBsm/OcR/IBoF5
c6zd53v7nTxLDXv9ZOjHjY0JqxtWjqdUVnyY+WdYErqop0M5+74g1LxXSBaD24qY6BsgWVqn0286
u/8nxLryLmmc3mWWqkE5nNaYr/9abMIvNu0bvNuSR/V9/47Gb0gP94ktKby+mIV9HqeUyXFHNxEC
9CDPHdPZ1fgDZe5iBFzhHYxyexFHynO974txc1uBpRxTlNKV2d6yNxfHiYQ7Mz1etdfEMSrdAr4E
BsNIC0LQ5hQUo6SMS0Vb8xGUckfBxLxpemMX5y5JuYsgm06IQiqo/6AfK04nDpFJzeyVjXUb4h2D
0NOMMNhP0jt1z8ZBDAQ010vek1eHsr5GHHJoMKqIL29gh+av2HuJmuFTmLpLSUrjL/WFzilZjf/t
Fbzu0K3UhOjHdtTYX4Qh69Wkn8BNGysNvJgIDKZMcZyqzUGc5ehOrkqAncwpW3quUS1GuxfLhcoi
O2G5lqXMP9mFiRI2hNFHzUTK6Xp1B7RLrTCZV/9HqHYvX0FnXgjBq31a3Zz6tLk0cHiqHrlAoxN6
XRizshYKRgfrUytUt3YcR0HlZGs0FPbFG9GlgxKfWF0zM0xH758iQg8YNpe5jxJ7PJ4YkfFAmnF0
Egz7S3p0WH8HrPMDnQiRGNYW2vFtzjHa4/gW+O0/VAEcPCzfEO32CFiRuuq6AbFE9IV7X2L+7Uc+
sbcAEklFGdlMb2GAz4ayfQE5tQzXIq3LIP4nV2Jx/6/+kHWqI4KqkFX5YSOAyarKlnr8OaT25ROs
Dj4C+Mpt+DNi7JwJitDGN2dmdRVASGyiN5UDigflSW5MvK7944DQ1g8vCwekGqFKrK+mJk9eZ4ty
uNdkt9N3uYWdLK1d3pfeUCBnFVX6SwOclSguKDG2q8NWtT6NoNCE9mbxGF9Y39IV4ldRvYpPWX1M
Fk1uhKELWkFeFqSLRhzjbAEAF/iazIadyMcxU3q0sca10qb1MVw9Qa0eEpld1Bg+jgaws6999jXP
jTELxZwXevJ/HpY9egsQGwpy8VLkdVs+v/OGZgk2zvFaG22kI9l+UTJGXEwI/AfSlaih/nFpkXN5
FYQJ3uqna9B+zu0BF8TAkdA1Td3FOnAT6SY7YXuXsPEUyqYr58/BCmN7r4twCOt7XTv+3mNj9L5C
1ZYXoftgesxwdcL6jtievulKybTmzlPyTtDce4dVNGn54xriPWcX0jjSJMl5r53BAbbZp3OAz0TA
oDIBGDealx6JNN1X+rQqYiVb1VEyM3dNBi2X9LEV45MqAO9F7V+l4vLDz7DEAVqh14rZpBz95BU1
ijqSJjDNREd4D+ah/iSTZ2WTUn3RowoQBUvx6lKbzrenzuIiU3apQhAkyDLminTHjhHVQhyPXLeS
Rm59hBXG2K2g1UdwV3Ss1STLEfIwB50gPt7lNkQAJh8PVHPlAs+U7xzxBU0P3KQBYsLUDJLXdDxY
6QOw6Uukd/qMPQDid2nKZKP5aVHVtnJEZBHAWA5Nog66KytNgZQkGbjLncB+Bh0lvXSk/lM7OSBl
tD8ytin7eSCjEQsiR5xIkjpnn6tahJ0RUiukCv+WbfVsLLPAx1nzgUHUn1S+jNQJZLlhTi6DjR3I
P1+TGZdpgOnrQhBkkCXRnCuCBAIOP5ETG0sqPAcIFH8JcdmpqyIiYo8Njm9KfVaDFZG/zWzpK8zE
RaluBreRM2hgjGeH+mWNyt+ZetGnJurnxTKT1JJdySTuWeuQf23rjERAHASwXV0mDNWD8ykRYCyE
lQFui2jVtSTWiFweqONWnLjCdaIcl0QtCO9bxGLKEsIKcYfS+u2XXCV/OY6ZRKvmQjLZdjUHZl3e
a/62GBTW4SkK47rtdi5K/VkpkChDwAlBj4Fj/4LWAnFQPtlk7a8sZ0JC8RqLEEAFiHtf+WHjChMi
5zAd3tRqAQH0rtJ3ws0gkTlbCx7/yZoffqUCyHgkBMresEj27rrBsj2Tmk1xQPsXjBAA8i6E343z
d2W+R49VeVTebKqlsKDXnX9DyXkaLJOil6714r/h4zI9q7c8o4jWz8Gl5Asn4q6FMLAiVAA8ZVml
S7lb+NMm7XP/P15G1v1tN2J+Ew/vj2p6bD4rTtBPUwwo/0Txj2C+l5a6c7Zrc69Js3K22bsA3Kfe
S8eNGBdc0rTZonI1AtsHUQSrc6Mq3KNf22zmfDgjgOSjiPyBFzceo1mHp+nZHMcogxO6TIGDvgqu
zKcEoAqprpfn7Je0XqJ4GcLPUKyhT9ZpPggQCfUKPGz6j4DIhfd5IV2FyLF42bstXT+e1XrZ8bQR
5xRVioDWImfNIcvuPYezByFfIL42iEhzQddJ6rPjTy/7yqGW1bsbkYrlYCKhkxh6pjmDAP4V/r/9
Bf8LkVyDkr0FN2FYCSBwtUuyz9c3XbnZ1towZQvWJCrXNtUBAvJf9pwbivqIc3UyZ7rfn366nPdP
RWJqewuDCvMxCbX/K8mLc3OhJXiFGn82BcExTERz1Jkc4DUkCkIyVCJPzv1CnjNasUnJxKUNTKKI
Fm+sp6/0cNgkcG/foPVger1vI+NyllpkKjZg66qAC322MqaB4tB+33SK4dZS3cCoKgEVr6uLoDNU
kkRb31uluoA3S/MPfd+dAaCVRXnTaDB8RK/oXrZ4OUoD6fNueJLXdPuGg7x+FKomv5wrOAztYCjM
+72GkB7R761qp+aqGI4H3H3+2k8/XLKytCAoWYmmpEHalySHP/OZvggo7fq6KPQz7DsWJYnlRTaK
SsRveMwz8GfvF3dBtMc3zHNptCtvnXWxXHXAi7toK5TUpkFMkGlcTTjJsqrpBCpfjkqn1Zmok8P0
lHR1LGURds2nai+zwaQBGYbVYryTFFy1rYgCi9SPJgmdgHj0uGid/nSv5J8Ftj47KHCkAVOp/Ae+
PhSupUJn9rsWVlzKmHWXjFDX+7v5YPOBPrYNi5BVQ4Q9MwhsBmetXRHkR6Tjs381RMxHTcyUfUGg
xkMPDsabOQjcAXoEzezgTEa8RZOjD1Lp73SEYT+6rD9JR3Us3MEqH35dQ6+QH/KzVRBwdt8zHaPy
tB3LYKzxEdBCk9tmMty1JMRiA6b5zUCdIyi2oeqdqrsNxsGAPZh4d2ObVgHEuvZYThnlb8A4W+w0
Jn7YFzfqv9wU1F2gQUzi+eXXusqy8+pNflSAzWYMIekxEBn3ABCHHuJLxMoZZxpLXaOnJhqr18XW
b5YFLsgE1zwdKZopE3K6aYoILHQLefDxa1cquOFvxpYzr3XWCkBuIwim7j3/xRIOMV99Bop9gcGz
SUX8paOJ3o7TMDbEeKT1+SHe7Q+CPAAoO7NxXmhBWzcM0YuCiaX/b2cnekz/ny6sdexLUmP8+lGb
5ndBKdRLlc9Y8uTEUVWtSTEs7J3M2rYePQXWkWAOgqcu5mca/Ehjxgc0UB7DMyDMJ/1LweCCxpw7
d3fXT+1Iag5KujlbeZ1qzSX0wmHP4Lowcp49JN5Wb1HULofIzBj6o67wPkvrs7aTNIKgyO7B6k1H
+TwUV7OQV146dRTUAxm/2yPbhl963yoawS0Kkl6HuFYRqfKTkRkvJtYNaNwPbwFXKqVM1jqT/Wpm
ezv+TcHE9QMIj7gkidLd8kRLv9GRXP+Yvqp838Og1CvgiVULfvS6WRPiH92l5tLvf7SboH2MEQJt
OLV1oKgPQ08UaZ+ijgVlL08hwTcBUslzgnNYFAAcEcxjsYFreu8CmieVQHiVWCQZr9tHir/b+9x+
DHn8Vv7nmHXZnbOPl6vboueyh1gxwuJyzeA1eHOt1IPwv8gD0r24C8+MzcNS1UzSKEgatGDs99j3
Bs+lIK7KrvkhL/sioS8yIgV1filidEuQP9j+P9BD05z6EG08XyJoaOIFwH1lHnD+GSZ04dqCrS6/
oKPVdLHzNzgIpdx/qatVzo1EVVTTpNCsH5QwKlglceNsNxK8YgIiWS9/XBYtQNmWxh+LvW7iGUbB
4mFgQekXq3OHsUomL+fb+VDYZT85xFNBR34pps0Zo28+rTTSoHw5SVj5JZZqgJRtuBzm58CH2IMU
j1G2Wa19BcxSvVJm6xT/pmPw2Jl8NNSrDkSBedY5E3k5ZGt7coteVLCq83jpBa7LW7IS8QohseVH
rhvkEqaYOika2LPdu2Y/v1ZuMDGiCMm7JKUC3zknuuD4EM0LA3FopNkwlo/M7elL4eibaZbsBP0J
I6AV+uKzD4wKJNrrffHwdqQ0+Tq12894S8wfTUJJD98Pz9eSEy4puWv8epTa6p1ugPPclxQbwUIf
FIsuGGyVDayQSfEggICgzZAAb/a0VYJ8tmIuQt3YM/xOM5vxMMG2wmJCR+2Q29CH0GAA67iTyhI6
Vzm7CxShblfDu1u/7ZxxJutJputgtHXHcNuY4TA+CGqgbT9P6t52w0uqrIJMLmrlJQltvjjqRbv6
kq2x5ewX8P2iKXSlflKY7Phh5ilo7CO8tISHEzR70R9l1goF98IF4je3eOLafjKaeSnThX590tKc
vytilUmBL+U/1L3QL1qwJgnNS7bnK1t7pUzTP/TP/qCI2BD1PPstL8Ngv1VRqVvg4c+0QRBXT/0l
qMCb+VC4Pa/ZUNjlKhY6/mtfz2/mDstVeodGxiEi4P0ZUfvHkRk82JbGa031q4J/5av7TMsmTwHz
bj9OuXdxXNHy9wzdLoBFtQwbb2M+koo1giTvCHDdGbjC2BayIafPPJ6UZBX8oB7K4b1CHh/N27GC
K+1v/+p/tVuQ5YnnLMVd4F8SA5mTpFU8KqynMaResVWmPFqUA885Nyk1FtnCsXEkZNtAQ5hmMQZE
o+V1hzDXLqd9RSKdQHwdF0+aQnCxEfYs1h7J5HMFvmdMKYqmLAUCUiJyxSKYWuf8988rZcRONslp
Je9eKU8+DPW5C8iHvo2ztKHKYlZjFlhvZRFd6y7NV7RUGK48ePx3zsgKg2vDC4GUi57InvGmPj3w
RvnSwIQLKQS41MEEHxeXgKpkpf1Naifa7tHJWY9hPu/U/M/Nekc9MbU8eB5lW8Ugt4X74+EuWrjp
fm55KY+ZQ5dIQmzbStT6DOLSVGKa4NBv0rC62qxsOdg8AEN328khKbKkZEyrA3iwd5pSCo65/daD
sGyim0rMP8bzDYls9r6tBxAafcMGp1r7RZ0ynrgdYVyKwM38O9r7sVTMzDFXY/DjgIizFRfj2SRT
9Byvx5gnIB+uw8FHzVS1MaZZbRPaDhzkVWQbcm9Kirsny3q2CRknrJorFtCDzpSidGKKeW35VEZC
OKoqrHwhCJoq7BV3VEy49SzVoEl1sVQneX0Z1/nXEXcs9H1f718xb8ApkZAwsTtumexma9zoSDtE
IVqIJaWgr1DIP2Y27E9H/vWfV+E7JW+JN5TUAnO3p5XBjBbR1p/tH7ld/W3ZW6RZ4bPrfDPGTKrn
ronlE5DkMYCuUXw1Z1+eO+38XAd1D4es1dqu5Vwop4ochzCmHW2OF4wnt+F7KafmILtMfblsKitJ
v4xd6K4F54WZVPv0egU7JWXAIMsWbHeyGxHSjs5rDkeIuhewHSMCk6dHHbaTI8v1Hc8gMsNeIf1G
UZQxa+febj4Dn29ktlAUq0ucqTMUiPIVpa4pRa8ZRkMwvGP590kSj1deT0+DMsXvSByKeFqpbxGx
hgOPS0F22gPlpI+fS+Qj7HIVqJsyX8JtysDHgTAvO/VmH3/5GiAZ2sKY++bgQyskl16bWIY+GqnN
WVD1PEsGDo3Bsno7iJV4Q6nAZuFRcaniWbl1uSyGHJSgLerVPv8ZxPfuAXK30/K/KHRZIfqyWYNr
wQdm3eSRmEGFRRCS1+TKOPZmZMFnpq/X7BCA578ZlYeAG0RpiiwYmj8d8BoxrXkwWeLz3bBUfNFF
7E2kTyDe1Vis7S8n6GEUeMKx3y9DhugiIfhHd7HFch8/wyrI8J8wNzsMHC44FFB1Qxqzfm9MCjX8
IRLKWnXAJlRIWu6UneDR3AhBzVGV7M7OU4P4TXhlPQKHd9MTTQi2zfUhGzi4jofx9CNEAfB9vsXi
pU0T6jlxRzquTG6iuvms5BvljhXGN3ZIupUnVs/TS/GlrTqtY9yeYxrOx3Lh/vy4zd1708xv6xM1
tr2ct/ZUhmFgu+dds9cA7cE/F+Blf4uw20KoWT7mo1a8Wy2PQ7HLH2iNbvajnX6JqG4AEMkcwzAp
zZssSu1QaPpLYHoCtm9r61/GB8Oo684FNe2r2oBX66fpA+0ch856cTSHYfEAL8cympuiXtai+5EZ
fwms9cfpeQlhfEH4WmezN9h/PWCUByUUsIorFZ7dsEwiZBF/DVYb0z8knsJ8JdgqhxjB+2W1OFfE
lFiHvyXnR+rZYHa5MuWkpsHSUezg+p8wJQ00t/zEzopw+lIR/lL058HUKSsZBdjWeIrnu8JVALYb
g7wjyGZzdsNfl6jiwcWW9eE7SLuLwF0gNwlZngSMJTEf9qwlRkRh8TKCSzUbC1xV9Nk9MmhjAFBz
FUl0ZqvcLCs6sVOVwrKsdx7KcBu9/SA1ngzrJXbg7iKpepdrG/d2Q26rsHXOcbyhFow1BNkeTVvB
dLTDYDG6e8oK3Gnm0mku/EuYsMhsrCZjeLSJZ0HJEMd6/kQjjIptnqTqygovmH3oC4dAgjx5GM0I
6oLmxYCva213hhG0Q7DrqIYxQ/OzckfYGmNn7LkPa64tWcG5z+TfagcEryeDcutc5DJCi79kDKrS
zjbXahvRIYazFZxqI9p6EOvcdFciOTC8ja7lxUMozNn3GcCcAclmmuQUXUclqZ5Za9YQATf7x1ff
s6XtDXzvey8qEXGbzEx5pcnwtifrKQB/B7vdi7uMgpLz10Er3hKguYU7tQ9gBfHi2y0J8eaxvWiY
zmkF99PmTNpm/RdovyalkCx8yIiFXC9bFjGbG9/C4zcnvikWnK01Jh2npC/E4wzkC83sej/5E5Ro
lGsmtrQOsbSlzDnvJsJS5azl7fFLvs/FLXnGoAcJ5ry9nsSwSNUVMUErDl2JMgRW7UDCsWxYbpNs
FOF0aqm6HbhtFQR/cUseqmCNl81Ko+bgv8YP2LwRyXg2NZIeewupoqr7INiyMQJS9F4zKHHhM0Xl
QUta4TxkS/zfha28hN/6ILxWIzSR4TbuYUDQrVHTL8ww1hdxWHG5oRy1c6WN/BwAoNMZJS2ikLzx
//0mVgvUqKvc9TMFWKq0XJqaG1qdzmGHiLgsS7WFL+SRtT9t92SFmWg8s51R+FFEXO07fHxPOa6p
T7PPMpYSpT+V9Fnc06YKJVx9N4ODqIirGwGP1YfmfzkaRXl1uivl1X+0P7xXkRaHaKN0ifkJvUWw
J2bcLr2AVeACfON3Nvp5Ac7WtUKYbaxpblC9Vjlc8KgeTMCrR1fGZ9Gv1egMW3seQA8ecZRTyQyb
3jBYii6tIa7M8uAeFXiKBg4dVGVg5ap/8L5oUpeRgP5kdO9HVrQTAKSrUYEKGZMZCtqHC3mYxhA9
d/x2wUVfr3s4DhmxjZwHWJdKlClxwCLm3R2AMl8hgLT2wJbccbl7lrzGCuFrYyZMkc8KYbGjQPVn
Wd3lU1/Xpv4zmwyhmnoyLIXE0ZzOdvA4bXjkgNpsli1maq1yyP4axf1dcsYaYgOJxa//rSJ4nae2
56jOYT2LXyc/izLz08uVADF4F1yW00TuuWTNAWueL+YpNUvn6S0MAZD019ktWMk0EXNjmumzZIR0
fQr9NlvB/2rqtHR8p8rlJVGT5D6IWGgRo9h+VVUPRfhd/SZQntL+BADHZ55zhh64IWgmZU1LjzFh
lTBV1yHlWbxE3owA4oBoe9ecpjwWHSsVb6pQQaipWbup52LArjl7UZkQTP0ChgW2Ua8ZTnqOcZIv
cqUEX73F5b3FqkudMJwdvRSvaU9OWX48S62HGCT69Qc+yUC0prxGx4iGJVwy7HSbPNJD9XiHM9si
tvP9qH3Fr+BJssUI1epz8MaHixU0j0xxg7Om9q824NEj/IuRg086ZVVryJlnnkSG1igZAbzIb0vz
5TeEhIAJudarNz0j+J/kE20FMnZ6sdX+Ll8PvNA2vC5EvcNuvM2Z/ZUNjpnDb5k08fqONlbP4faP
4+EZwhn4YM9nPu1hO1nWaa/itdiBYOsKnsAV3LGFSEeOenz/Y/AE8Jku/+KZrPbb+EZtYtSfQbXl
+eJFv/1V1F8khzaZva3H/vMdCkJQe+qIjDaUnYV1rG6SuU2lBdvBnVmtygPBQ3CTN0qkMvk7viSQ
aY9kSfNxRPi9i/HkgKm3KmXttSEncMX2J2TpBIL4Et1IqPxsIttT56s1LaE7YVo/SrlhnPX2y65C
dIG/vd78fV5oMgjH2M51ceHVoPbVEuaPmQBmyvMAnreNp+g96PFmSvyN7DOur4lQ/5IKbvFhDsCT
9YuYeHhZJy9li2E9Q4vthjB8klQ1EGHSdzA33YGXP87BFsXmabQwfF2x7PHWqSu04QGRWHzzKT00
Uj8ktXCz4TkRBxTV0VXhVjU7hKGmZtFd9THUT01JhsBaUm6Wbh90qoOpI3TkPZz9aptKRWslCUsQ
gyRg98FND/+7Jl0VOW8rIBV/eIew/p5+6t/WwzcwDgqTG12K2ysUWlLQNrKCR8FckqgNpG9iVZXa
/VFZ4yM190M1M1/AHfmBwN/8ofNMUWcOnTfxeaNpwOAlHKVPorNRbvORsrH+Txek1ufYv6HG38De
O6V9AO9yWTBvcZCmYpWcapMP8bHMqaUhKMcngIEgEPFuP1/NFYwZEGWcIpK3zGxfNK0w+Jm1qxMc
wRG8miJXUigJfvYML4DA0gai+xYXVEM9LaeFlQEWBqTJh20MW9sgtxsyyDH97aJXJNb3GvUF81qq
+DlzMhi+/5anoJ7aU2YklK00JWmmcfM1RUTigSkZfJ6iThfbBc7PbrX4svjiExi+EJQ7jQZqBRc2
VOaFjJxiZelAyFNLnTF1XOuKhoMZ3S73lGepPI+MsawBbb08bC7DVnMnTCNLr0c2hdrFHYpbt98C
5Mlc3FAE4zsqdK2/tFfYsQLhsSjVXspfDfSGmbeXZlHBfO/DseFjhjbTQ1TmT1dWgMoO6bvrDUtz
imjVy4a+RJ5uDsyshsOec+QWTZ3AR79CrNzxANtEb3XH2kwwI4HsSjk7qRsQvZOT0ibrRzSv5ubv
mF5lCtVIV57TN8jecb39yGud8d7I0gRuzDGf+aUEG8vi3QidkMsU/Al27jCd01GMHGWRklUnAIiV
jw3m74VA0thYHqIMpAlJ7sP10tCs8N2Q0WRNscMuODHDmK/ct301UiWO8BpIKjtUVb7uPJ8kVhzP
hqMCPrzk6wMMgjEvBpUsv166ksKWnrC/nvrWhB3g2cmtmpzccC49QWLBeNsQhkrari7yugjIP5JL
PVFWe86j1KkOabP39PYpKBQvsKXjZOz+yzUAViXWHzSaxXFhSlXhZrZdpFwVdu1TD+SrrCEdT46U
yjBtxisrhNW3+/aqilomSab8N6k2LAtB2fY2DWPpxXFi4M8F01R6fzK7R4DLkq0l/Dpj7PVJLlw8
1qAKXvisSFqG7bhKicejnXzCaDnBaCSZ3YC2lScse+UCU97Z09GVaGPfm7WnMnpeBxrKjROARZ/S
Z9d1HoWuCIaJ8Kvg//ErYZVfsLUIcdExLecHKfPM5ayvGJ/SPfQH+znVGFPUsvphH6HBlHQI9xnu
RvIUIVizohaGC9igNMFKXxaFeWKvdrmmMcmVjJvDjMAtxcTncFYK7rfHi+OFH+1yFZaukcadji10
sA3NP4oR2EJWIC55GpytWDaht6yoxsf+uCWV6aJTO2lMtts6Nl5gMrglcynI1l9uXX9sc6TAmInb
JzV+PHL3NghE+gZbfL3VvW48KBcSVQBghbjIhHBbYedErys7FjgnxooXIJ6wbE6uuo0D3xLnzIIu
09cAJIcjzDlKPGzj85UoMCZlovo2VuBflI5Bo2cTUEmKrMvN2ygcuRtWoOaeufwVQ3TM6HyAoY+T
gRiZblmI/qCYgOMP3ble7W0XptQpQ7ZPmE9T6+Y6x4a9LJu4fM8GU/CHM0RJ0aN0yqswMBar3/ua
K8QIA9p0RV5A4xWQRwQaHn0pTBUoITB9vnB/gQnYX6z0/HtPnA0RBCvjoYmrSSPa8KYsq7Ul7zfs
qJJp4fMIILpda42JUsAuiyODYPexv4hFtDv6wLCHxbY0BQk7BfxAKeQKwxPmsA7rx9Q2xgHaVodX
OK+PPqJoxETjhu0ONCEaDltabl1J1Si/Mj4w1AfZcbv/QBKcJ5l98eIgbmFiA0LuAoj+Gfwe6k0I
9fvP6uy62rlmLDkLiXvWK13alwO+/2QkSfz6OGZYVNgMIe90dx4N8Vlm1dJ7Ri2wJB+HnYyRLaq6
U7mquVWLjzGqmiEaE1lXeGrvSbUYsgK9qWmnb2bN3fEWCSQ5COHNRSK8yIcgt1xl96k/y25iNZ/Q
eFdWLHtfcj+6d0Gg4yotmoFANp+szdKXzBkY4JvNmS6lmUbrfPbXuK0KjyYogjbzheV1xpHW7k0L
y7N2IB8uFNpiw+tvIF313kZKRGsGjmwiijJdlgwcNou/12oNgHScTuOCvLoV2xeMQ+Xw6T/YwGoT
i2JSdxRWhcG45lXDmFRcEq1BhpankRbGpmM3pGPeI5kdU7v06N4gHwR372DHRyo1R/xWR8nX8CCg
FTfIllmWWmzidIRZy5jnWA3KHeuvcZ6Ga3+QP85s1sTnElMK0RVzXhXukUjYA9248BuQA+REyePe
kWFywbIhQysC4SWVTTumEBrV47HBAjF05V5jCcwF3UAKxW/qYonvTH+qIPR6qQVnRQxRgTJSidQ7
gj8u+lWr7Kct3z97xP9y0M1djAuq4yi/ludGFBQhIbj3K1UppYzsvlh42BP1v5SWr5mc2j6DW6Ql
NZHZFvKb6o6TzG5rBjE7AyVmWNmqCFWUHMC/LzeoDVSNa8edJbsu9Ty1narHhBmzzQDaHh1BXqdH
xdM6d7KITyVX8yGcq2XJxkB8XJ/jVDRMMd4czDhnXV7XVGTMCoIn63XWTFgQcQ+QeOQnewcxboMS
ltWnmvPXOLGPQ5tUeRedxgn+TLqdzGNI3k5Nmoi3v+a3w3ZMzbWpVJ4bCnGaBsxJ08+Ewl1biwaC
aQ20N3MzT7ysdnkimZdsrlIe1Re3ahhHyTMgTWbZ5XPhQC6VdGeDgwpLz3q6IWxC8rxDLtsLHOHt
voyK06I9YZZ6axsVZN92QNtnxK3bFiSZcaJANEKoP59w3C3flf7vZcZi+phuDK+hkyQrsmZL/s3u
N2imWwZjkNKezJRLtrpB0is+50nxr9tBnsFrQfVQ+oE3TQIrOtWzmmXyupmcGqMjfA78jrU9DYtg
R5fDyqHX5ANYLPQYaSjWg0Qc3P7he3sg3hMR8y/mShZVmF32TV+RiCHhhpKrMwZXFVnhvrK1Jeu/
MfiCGG8SZackTG+0KnuuSrM7SiKMW0i2MI1IydiRTXQa7uEaJ10hcf318g9g2b8KaB+zBBPoBO2M
o//pqvyXAd23g1S6YgCrEVbuVRyldz2dgOFXoMH44xEMvtBXU8NleA3/Znkd2b19ZsZNZ0W44aEB
IPFjja22o8vR9dY2QqtSNnEMt+hvMEsTB1rIbQcqbvA/MEBw9OmqsNfXt7p9shKXqJ5fPaGAmgLs
OGS/djOMgyuBM4d4KKU8AwrTEStXftN6a7IHH+k4ZN13LrbfS23xWf2zulgxzaU8U9S18nay77Wt
VIi5V8yrwx4XS7rsL6NWIlGWyzx4rEETg6X7MpuQ94XYLJMhJCT8ev5OZ0vkeKA8Z+YWzuRXM8zy
WVkA/Ai+DBmTqaLHqAFYs7fabh7NNRB9ho3u0THYsBZ6lo4vf/pDWo0V8tsg6u/8yz5fIOo4Acec
/1h2DjZVVjUFn+WAckyB7KDgtwK6q4q5eH3+dDC4FVgKH7IqE6tR9awsYSnOSjImEncoI+pwej4X
nN7Wr64SpQXtB1FyZkyvucgK+Cf6t+tdCOblmITy9vWXa2/FyRhnfCsFq73ntKPvzjeL8SpBgb59
mrodSk4sF0d2urqj4U4SiotuVgSW+462byGYwmm6gDZnO1yfzAhJGXUWlc9zJCG27ps+ForhHq/M
fTwn1ja2Dz8o4EaJZOf01jROkOI18iStU1i1wT9v7PFE3bucAXJXgMn/KJdSNG2I9SVlaNw4p33t
xAYXLBwKt0Z5rCQ8nQczBd3Am058X01XiKma44BISzVlppEG1Rjnn0B0I7vn6U7g20AjptQnO5eX
+oJgJXgQ2pdYFG/i/Cxf+tuLahL6PJzgB2dB5v+zdRR5fRuBTSCJpZF3zf28UL2nxeZQUpUwuh+Z
n7Ohfpo7I8fDA12ui4vqtlQ9Dfbv0b5PcryOPeUeaSxqvuDqlzywC6N6nSMuLYgj82t6IFlnY3/W
SPCC4MPlBhafyn/EfDeP9FRtUXQKbh/WUD2yWxPu+FZvlpgz2+3Bewli4yTE32nrlqRPgk0rfmY2
RUuJ7yuSbi9817HLX+nc4A5gLYf7xRcaOOQceeniLLsevCRozcLesLcSvTmfk4r0g4m/jCYGOSJP
q5N2o5AQblRcQGKwEOgq6qi2IEE/mgHiP81RPiRkPMfYZOTO4emKkN+qCGIfHJhHll5Fo98kjzZ0
CrwsbXF1VtJ9YK4T/ay8fAG/3Cr+VL3NOGZQi4uRBdJ2gC8yLzjUUf9MPhkMVthxDuscr3B0R5y+
7ZGY1zkXSOsxizq60H4fDo/O+WqWwpTKYKHLTrp9qz8qro8FVhYYNkgn1AwRftMA9Fpq2BFLd5aI
NLHS5E6nw5p5jl5JdP4RstTdQv/lU10uLAhR4cYD1b+yCYWtMJFgFhSrh8pBA6vrrRBSDzIwV8Yz
0+DklmxzfbpKI5UgRQeQTHa+/3cmoiOk/EXO9KuJFITvqN4389b+0aT3ydvXiD6O1KyhRrtinITI
/M+YXW99kba1p7pNx00q4NDRS1x0gZUbiqQx6LI+cB11T7kCdoVFIYI1wq+Fop+ycWCw3tmHo6f8
JwikZGGYi/WkxMdy/ilTVC5tkudmVL8ZGzLteCYIdXqBc6NxKtrEJW6VTq83W1mHZneFFHWV0t00
WD8W0kREeBcEskTxF8O/ddA/u2q5zbTu5Uu64UMn6lg2KIgtMo/geYv4lc3kStKXYqXOoDX9gtMn
XFn4/FDLFufXoT7urOcHoIgfTj2tOFPBSRVDNavcw60Q3lqGud1Tv72sT1t6Xg+2/q2x9Y9Oh6wN
GVkApJvS9YPZIOEyR4YCIoj8s/F5hMwdPY8k2pKTEAHsctD0tNlIj+P8IFNJN4LZSPVjLdlPp3bt
fmwqpIgn/MudeXiyQY7MW1Qu95vMJtxHN3P8gTftiU1p0hqttRgCck6DaE6VUc867dcnuTqnOPLL
1qPf4R/jrVcRsNB5M3hGh3zSH2FbVn/OPlS/jZbOvPbHrN0iQJiMF5Q7nxLEqd74uB/zecmAq2iD
xkDReW3xxn9qvOIVVWtu2uy6rU+eNvfkbfCyKBP/zREzg8YeJ6XfgWPFo8qkRGuuo44FgMVdzNxo
48Bz2Y5V6QGL4CTPTwCBSQnPaTG927XijB4tNS2MmFRLIMzuae7BTXNF8BMW3KYJ45Y0Pog5XZmc
c4fcg3Yq32eyeI+8DiIfOgCnkVXQds99gCkOV6z7sYX7QNG9hYwFCKIxjEDUEf/SEUnK1Ny6JQMn
cfzC9NV9pC3u3BSjFFrROf8a9C0LrbnLYdGWbUkTBi2OtIAJDiY35hobOcBJT4+TGAzuICaIrIeb
4t4vXMUkrZj/ABi3VX8XxlCq/rpJITzvNFozEvskHfBy342nV/3/jjvokCz5/ynbX9w+3XMeIV7R
pQ9D4ipYeXXvv5oHD3M+WF+UMqmJeaqcX0vIfDurLFIkdaZshnsVGeI/6OW2Yuktg7iDCYo6kQOq
jE+jXgxE2q5gMBAXz16to5yDgH1vb84QIRoWGa244rW4VbcDp3UuhidpPeqRWZBajRWuK4roEBWA
vjwfmVAwppR3dP2lME3qPxwDQ419VfwzXk7emlkXVtTPvXiz5VOFA3lhFVyOO4Daopvggw7ELMYm
YUGSznFRRE5+lExwHPftDXGMUGXyshP/PVJM2tqvG1pPdgVWTNM++H01V7DN9fR2WqH0Fmod8xMv
SIrAsWrvQ1ehTfrrhAdMfwLH0nuf5e683nYRaVxGtEe1eYEBkHvGyyILcUP0rNnKGYqgax3U303I
OGqL+ESGFsKZC3f9R/jpopkHoXPOuF15VT4D6HCFnZElfGtPLc51iej/IvWqTpj6JvHDpFr6seul
pQVlEz2cDK5JUadZlJfSkXT0TN1hOlRiFuWwfu6TL12SA2+TKWhL5RJi/+tr2YAu9kfjfTTnU34b
mRR1np2nu+h3FIxFiRar46qBAL58DbWODRMz9OosBNiRMwnpKVWP6xdYkR23nQ35sa1+Vys7mW0h
MlgEpW1aymzBK6RxYT48Jbx9bncbSdQnal0s24g4RtFazTHk5/mYIDqgXG0yLRVf0ipTQWXEnqVD
lOeE782MT3Pp+WnI0NrYdlndEl0HXC9eqDIniPH9JhqbtMYUdQmqdqr9KgnH3iAyYXgtQ7Wtk2/3
iTHjD/3WV7eL+RCX/GoNLMGrT2+5DvmvAYvUUfcS12lAZfbeW5oi5TX0uXlKfrOwlOQqpfXLZ7cX
ZMKpdy3KVe3ey0CgHtya1Mb49js4zbc5W4u82dT+S5IrD0khx37wAkLF70rOSZZjpey9518YFqPF
3rADOyhRsTwnTas02bVWohf76U69t7ExaPzDxVc7ogP4jiJr2GUm9iP/6StWOPqgXx9eWXxDjnfn
tkSKnU+LI5EJQQQKMlz77bjhiKAlgI6MB8IPEnlnc1lGnbMsMPjX4Dyxwz0qqcaEGmxzySodvCX8
/0mzp3tc7tKXBEOzZH8Lv/Dub5R1Wq4rXL6j69IFVtn0IZcn2XxkwtbVdC/q6gxuHTNs5CYNiitc
FqRh8WAZ83JB7PEqtIzHwJsYfCvPkiMhom96KzRrFeQz8+mH7vtAo0hwRtdAcdYdvDona4fBFlV0
pv4xpSUNHlBFytwSfDaiZzvNKDovQX97S4VylJ72J9eGcPNSgweV4LJa98Tpe+Kyu5WvD20P2f4V
r0j3w5qyJ8qAszZs9kS82sw6s5LxpaAijdmAC5VBa+DEh8rfEgjr/yPNBnjTp/O7lep1xV6+ipaf
/rAp1FONSaamddtOoFnq4bt0sCpbWcb4+WC8B0AmjY80gSUT5cm3utoKzz8U3s7zFEhRJLEQJ+KY
ZGEkl2ShvYspCJHKf8UibLjQEr5rJUoM3Sk7IF7bWKVzkJcFuJ8Qnpwlo2h2DKiCfw01MfzUXYHR
HzDmP2LETny2IijD8pS5QFDwSkz8nrvzkEHVm5zag+aUAby5Cbv1Q6GY6ya3llLdVhgTIeivXKnh
6rLsjiQfwJrqM4n0tzxb7mYRPV17NHC/4+JzU6tJyvrdSVf2ZrxGvuCDSet4pMa7fGAbn66olSQs
pP2WD1UKeKDgUeHCcebmdZ1Ek8qzckYkktRCbLXlsS1ZyNhzyPGOUw8af0teMCBTsGKcLQYoWLKg
k1h5oOUAUP3oFt6ASB9Kz2kDeMGee3c+F8cyBYaG49MScAbMzFd0Skxk/9WlRSADX8brhXCzYmII
jRJRgYle3FRbdunyMt08gfEtgcBA4oo//lDjMHz3DIgJvJNspeVy9OrjWyDxWEVLSlGsqkfoyAHi
Mr4fpY4G76qyH936JLzGaYUGkx2Knp/X6Yl9AfMUx2/giTPiRTjyP1nZmM+iRuTDQhieAMXK8/Qi
3EQrUHgMBxCYa0nPHbo3P+2NFvJSkM1+dosi3yS2o5ZBxVRaOjHCPwz6Q2q2SBV6doXtfhJZ3iN+
Yiyp07vkTEPfzXs8NSEQY4GFWv3EVVoqpLC/JQwUgXwfTOrgHii/kf22oWHf9oHa6PhxcyMTJX3u
L2W02hB+6y00iXoLhaxhfDrKT5rVw7frhchHuAx3zqY4zBovRZZu1CUfv5JNLI0dQh6k1xbhOFum
Cpr47+LEPloi5fLwzMrWQxKjaFQmq58O+uBp3ABO50Hn6QUdK0BkTJgvpjleceiN2RGt0qO58EPu
DxMq7Ycs6Uxc5iOJlz+sbFZQCpxRkwznKDyusDXMzH75Izlzw04r8hIJfjIvDtI6caLJFbLS8kU+
jPLLRQ8YaG2lwQhMIbnXU6/UIsidK63V+H3Lp2Gz9qF+tgjBEWuWQDRDvZ+AMt32Mm16Vzbioctg
/Cifw7N3xERT4cIqLletEwc+H3/ENF6m5YuLfinEE282ZLlE/q8sqtaBhAukSdvFZJvBy/St55Kv
FVAw1U0T0o7dFln6TeT1Fr9dww3SLU67DULRWYAR2aOa0t96axvaJo49rc7wWdEOljueHnylTKcX
EwXTjUdLGQLqUf05xES7OZdszuI+bWvlH3MewXlNtv7gNfNpyzGYCEMRqjex2xyMfpdIQYgtUPWM
zA3FtK8OvggcBLAxYjWLT1shbCCmD/9w4d7KW/sRX8GP/HGkQ9D7reymZ2x05+X7e6jVO1aDd0Ln
3iQWpWLQFZdNcfvonpdWDyfpaU4QwdBky/Lz6JZSKQFSKCS3LY1ER0stTf1v6UXtdX6Awp1JE4h2
wOjF3PgRrDfdOQvIDdfOQfdMVCpTgxH8vDokOXnuSiPrhzL8zdiyFprnaUNUSKTsFIY8x6C/g3LR
QDn9m370xs1BPVnmhzuAP8gR6LJPY0zPG1gstezablqB89YFSJgvp18MaHi/4t7MtV9PgPQB0XqN
BOzslk23QtWN04leqryRSE4rbUservVFCDP5JgwGaZC3NCN2XPM5OtmZrY7JpiPFpYltnSbtUj7E
hgz7XnJcTaz3f35FH1SSsO/sShGFgZy5EbTuNlQU+byEi9/0kGWEViEynPS8vgUNpNpjUo59ITQp
pC5Pg+H3D5IcJfDVGNOGRA9ZmXmih2Sspxo2zjXdT/ShsPc2FX9WhjnIO5pn4/DH352nN1zvN3wf
xx0nfq9OXDG7LinzB0KNW6PaBjfZZb0egij/zUrvZL+MCLnV41qfoXR4kZfso4oLXJj9HTtEdE1h
vKr6RUbC89lAJQJbUVU/LCIAf7g4EMHnFho1wiSfGV60ymGrywWGkUwQpXEhyug6JMho5/3gf6KG
hrzFYOTo7UD/svfTaRD5xt1CP7CVJOKp7vNSMEbwT/Z7YLnkywUeWOtF0KXnOExaf776YBjaTU/f
GHRB9ugNvzuzjeYyUm3QAaMQO/svSzeypBrYpeJMXYBQDkpgNX5hYikT2yrn/quqeq5/gV08LYov
zBc9YCP+TjVkKI9EGcrKi0fvpCl2lyKglzlG04LB510iS+ywIB5rnuv5GPluk6hDmTcnQ0Jr1nDU
hgYEIw4txysZAaD6miW89vaYM5nepZWeVk4hW5LgVzDleyxKBCeDiwwhGFsNpuFMkcTQI0g5MknY
6zMd3k65Btj3phXaFUCzxoAEKPsBznORT3EKMKxGmoUSMGoxRdIBAWjtkRZRtB3DIqDG5ktAGz6I
JIuswYT2fT4lM323z1pnel412Gm4bgRsAy7c/TRFvVrQR64lAyW0EiJelpC8FD7+/WPzmav3xiTR
I/UnPO4NVFbS/c66z9gr8jVdp88DAJLRhiLWfpTjc0ZjYStKTYnEldl85ofxjA9RIdzIWJRggqm5
lka3qoG/wREFmUw7WqFmvgjUpRwhJsWEze1w5f9l9l9HAH5lwn4dJKVP/T3YIGLHz+DHDXssDvSs
15awZ330USsNq4MM7tB/QICgOZNiX1vuSoeOukA8Gg+2+J48ZG4DbWuKpL/b9ujt+020VwDklXaW
Tng30cM5nyIbUi++9HKtADVexJFk4ePPVVIzNvB7JyYr+XS/KIzqNzrLRgCBwhBlMZnbUdapm8+r
op2DBZij2rh3eVFW2rOmW+UlgfckDRK2c3a57TlSkNyZFMT+J3rcnQUI/3PszFqsTEB7AcZOOLmW
SyA80TgRCLqr05woPj8j/BPeCc7HTO2tRA6Z5vR1D8i3eh4eeGsIeHt6caTiGomNsxhH6Sz5LEOg
gnZtsccvMhDbphqggQf4YbtGoLQJ0cDrVY8YfNURf8AxdHY7uqUu79N/8mLK491KMDBmabKWySD6
IE1kHOUELSAjWnjN0zIBkfVaT2MbxrgBrBOVwlLPS2rwSxIDkekEK0NTpSGIMywQY08+FgV6BIjX
ECNMSaMaGg0RqYdEoecBuh/1ddxyVQZGHbUioWlS1Qp2ZBPJolyoQcfa7BnBZwC517cvot/9tYC1
RqCzE5zinv9KExyQ19JkVoJnXGDtL/3hbljGP2yBG4SEQgz9mT04z9U3M9sIQGg60xOTKwJNJFTs
LmQhfsxXAvloIM+Q+f5MIjR1wm/SRubwiwM1Nuq1ODu9eRTyfhp/tI+1c7pmdfsu4/lmpHYMfa3Q
fQClkSUnF0VZRj2lfeWwVtVKgZR/vkdfID+bynLCcN+35MoTjv4DYgRZ4O0h6vy4AJtAU2d3Wrz0
BlwXuYI+ROrtD2AlQ+CMvLKXxpkFjO3nW3mzmhU7swByDcywdq9yBs/YphgywPtodGt27RNpr2Mp
3sV0rEpSelTUCiJF4EoXEBP3JSMUwhug7wGFeVwbO82s+SnOWnZODO5QtuQvx2DHV0W83o68nP/E
oAJaPWp8E+5j2BOdVnIDka+FFHwDbDx2uFUmGXo08X+rL8KBck9aKFUHYmuu8I9NZvbAPX6BI+vW
CZQheg+JZpR2ZttcqlCY4/avgBkED3m3P6rMb0a/7vEm0FNjoHJoqUnJALePgyW7LZRXamwc80mJ
6Y3IYAFnNtgmzdcPdHogXCci5Im2CEdeReRXsR5k1aKgSdwMTfsLoL5mX69DH8xl2BC7u8XzAA4z
53Ps+uP7/vdIrMoy/v6eJV9bCdUlskhE7fLf/A5ZuZvGSmu6z6oyPuq1Ub9XhiifV7hkibGesmtl
G4jtl1X0Lgwj9DNMBJG+x/RpUyPUV1uct70XXweksaSxjPNxtSoFbWbmDpjtHjd2sCmRzYcXqF78
7uzIPQ9UuX0YwQlgjlrZj1Ijb8c2/If+xUrX06K5bXF1VN7s8wGjSMASuEIxMch5b1A9Cs479ofc
7sU7cxJJx2FYcKkL+2WfkQovZx3rOJkj3DNxLuxaPhEu7deSekeH7KrbX3wIacwRy/LvHY1+y2bt
Hs9G/1+SL0le3Crq4nZczXJuxhdRImXclEVEAFJmqgZJ18DTU2JZ/GZdtCUJoUJFe/tMAxbx55xP
TMllEQuglLd3nZAgbtEkmBnjBawqjEj35rbkW5nDziTmSXdcPDtU1eFKW8zg2d/DaOL7bGH63J1W
aHb10xS5e3UfE6vBWq4KrBPOFZm1Oc9CsZnU/2KEhTNv9eeVSFYWqB1t1J4BZdyfQrPCdLMIskto
a2KggHmsWncFWmJ6Ws2a77sTP4ec1XIDRZrwIIhmdDxfKKo05dsKt0ZNT01PHMdWTRq2UVVb+fyA
X48tiHJyrHQBs5+GtVlANvMeYqAj9b7flE4iTSpn+3gF+cgocgr5K6iNcYYaqwXAK1P7Xt7K7DoD
4vv87jgUsjRSPRqhEJXAeY88c2c12BUBRnPWsbHglQX5w8JAqDhpfJIafeaixwVn9wGF/pBlhdxG
fhmGSNQBno2I+UGUHunbjvoreEWweEtdRVJT8NMbi6TAz4g65bmBXUdL0mNLwH+EGY93W1QsVHLu
5AgQEzzbEhEaHRn9Gz/u23VLy1q1c0TDxDXZ7vS8o/s7ZGqpa8OVr6pm3yibKE0FRpZjUQz/arG0
kualcW8GpgSQPmOYyZqpWM8Nx6OJEOUliRBtFvh4DBqj/qsXTIevL5zv7CCtLFQgkMqkJv0/Tgwp
ByIqMtIKGuJax+RDPMOHPoPnoMi9LMmENzf5pyOmXRv/5yelraO0CPzmRsheWrjWb6j9z7pxTT3l
ehzn+eZ0Xrqdx9o0ByTuIdRwsqkidnzO8E2Y+Lt7hTIGM2mPk5MCa1PZ96DnevnqKhYzOoR1VXGY
50qv9AACpapfbn1wwhKmliXbgaC4qm6kwqVt19n8S5lCGrzvoCTmUIo1fLl5TSLD0znyFf/sibLh
dqivnLS2mv/zyOkSWVSlStjA0NCaJj6t61BbFSeUc5h66tS4U4AXS5SyPtM2ZwxG827jY3AtIJ9u
Jjqhea56o1EOtmkOHqa9JeNlCzINhl/I+aUx2JrNpdc9jUG7EnrUBesu7ptqcJYmmGB0MHOrRfZZ
vHYE+Q6OoGjum6Ak0VNtKM0h2msk5PFPaOrTxG6SL2L29dTVcGl4pcj6uaUluSKfwt1eryJ6jZwN
w8FKFGtP2ssJH4KRanc1z8040pCvhdveyWTXWIAT1UYAanq/3Z8uIIGV9Kh/PrV4dFoUyLgtRLjy
Os/QWGiNJmpCvkkyr6nHK3l1PkAsxvxrGHQq471Mp8LaTCfNZuWE4zcrRrwaKGqvsr3W5cCSLO6F
/WA0K4JOD49aKdIF3bE/rk+OCwbZ2zIHlDh+YfjfxYUuam3YotbqC1OOpy+qEGavRS0zEve9xQBY
D6CkKhZzq0yPYxUGrFj8bcPdqUC3tVgPQzYSSW2gHujx9Ga/QAaRfWpI1xiVRuwYoSKX4eLcvuIj
tJHQ5+yFOLgd5zJ33uwqfJKFEKv0n/r129f/d7vMS0I7R0F7EO9syKd/vunFlOQ4l7/BSZ3zfhKG
6EMhzlqe+ZUsH+QJRCYB4UyDEG6Q3949KWJE3/V6DmLMx96wGVHxfaxZopVpcAw5X8uWD4HdfnJ7
9J9Z8Dbxbq5SeY8gUJMXk5FpgBNleud5LYSQ9wgosoSnz0UZY+i22tCdZR2Dfqz4prHFMmp1JD9l
IPpedeUCbl6R+nV5+DJ+p1fsdrbB6O7vsm33V/m6ENH1/z7bRKjAzGxH1M66oVt4kPgqXZ3SMXgH
jTTODzijVqfKLNynHD/6/BAru8/eGa5M0zjlPBYMJYfKo+bpnOmZ/ZPRgGv5FDPU879H7NzX9hZx
YS+ry4dqqAQzopdthtu2zBBBqdfXfjEIQBzSdvgSqwkMvp+hMJQWALsWe1TDlYl0mM0F6kekue2D
FmW976UdYOlDEML4/iVpLDWKRTKg8sDc4FI4bv89VVhSaJj0UxL2YZYMXpUvN93PoXB9spPUWGHk
dieGnWZLYxUHuY62SWzjf9ZSUwPM/k5STdND12PAqeOBSVIc2I4883iAtHUDP3hZtlOB9XhZTc+c
mZQozZmoCDvPsEM2nR8Gq7nLFE5T8GlPGg6+GvDR1I7YODsy5SKW8nd7YV7u8XrJorio8r0mDhoo
x9gC9eiGy8C+YPy4JRBZaE56BowxRPy9RQl/Hz1EDdWrO3zyTLccSCN1nD2Uk+M0lHr6WBQLr6TU
YiyTw40+KMqQJECQ7Nfib8YCCuTLsCg9q2v3S/9QECN/G6JEAGC4RLrk1u61RZJfR/h7d4x6DFvs
KudZkmC8n1mt08vBqfrdItj2XhxejxhMU12Hw/yL3HLQCnJNOWwRWaEViCvPPgrKr0Ejex4zSAG3
p5fNA0KKixuoqy8ST3d8gYu0kif+aMEOcXnh/w0KAIRXCgMF3er9XpZKpPDvobgYGzDT2ZjLg4kb
mlcz2sIdkYm/Sp1NEHYFZkGcBqdLf5pWdMpSd4T7y7R8Q5icZSW4pDVEsTZGpZ4E1TUw95rpx3T3
ZnKDV/1Qh9SGR00SzEqzSBreUirqtxR8hmpNaJpkCW2RLCuHM5hXRl/BBQw6QCJIYEsxTd92qsAJ
lHsxQwZizYR13TiZTCkYIblJaQ3xYjhiH52Jp+DkaoGxzxFtKOXWwyUrR3KdwCLEw1O/Lb5lYcp8
WJ8SQ71YxQ0/02WzcgNgeDwUnUDK80Gk5ttcEUSjgJyLfnYCNAhHl6cUiSF3q8LcpiFDdkzjwc45
34pJXzkIzgNGGLCI9uC6GtmWO7lYIm6ZD5NZk1wtIVl/aN338VlmfvT0WoA2Tdpg16PNHrYks/HN
YpBGIBwcAtleQXISWGJqqZcjoMr19soY6HzdQBeQc17f9JFjAX8M/9+qyZRrnFeYY9BpmvQSQpTC
1yTg0lzBErjRBoFSd5lRYWzlqWGtCt2OEhFoq2iv1p/Yu0SS/f3oJpvQggo76aMkDfu6XzXKz5qc
ouS9mu+BOiRuc9kC9Uvd0yddFHLASe+SvyhAFKjf2Ppegjg+vy2gAX1Pyf5CZERnziYblmyJGbfX
8u2CwpUcZYg3OgIkhI6Q7ozD+tgub3YJ7oVi3Asp7695LdZjk6PqKEsLp3flgmqUqYKVozrRW+lh
aRzqjQVWMGCm4Zz1lHMZxmW6qqQHKDiC2x93S60bmwoAbd/Lm8YCI323vQHZ6HDD3IyVdXRIRNH7
3t2+wjwXfLqt8DzTW3fClNd/aOq+sk39MouHfk0LKlRTKCITpkj+IkBSDNI2tobIP6o7sxezrKqv
JpMMGVIW/2TMOdrzhd6iAhtzuJkohcT5jgyMjLIAbAd4+9zQijdThtIE4fz1/+rMqL75ZuSmQ6K/
ca9ijYeCRQdbiMnwArmMPzbg0aJ33xnqOLRWuBwBN6LR0YZxF6c565u/afzS9CHs867eFGKyvvnh
fwg7b0UDnHISJa02FoURY1/dLhuPb61OXFyCXyq5z7jiQfos/MyY8rBSgFAXfI2NC2zjSpHP+7ia
ngaXHg6R7yp6LTV5G6OKYW7wqxaXqnQBkv4eDVrYP5CKkEgfG9vwnHTj93gLr7Akv5i/b7cW+tyf
zHMmZWZjKhBHeHuwODPPGZPl3/l7zV6fnTIJGFNpTHB5JNaSi0L8PVF4eWMUB6ew3zUoU7MZ1nI+
HRI3g84WN+152vKnslnO4iK7RBtP8kL5vcCECXkkDLzaiwZnlzNU+EvmPbi6oC3YtUzINF0PSmcq
3KxqeCyIkAoTwYZdwK7QgSK12kZZ4VhfZo1O9DVf/KcuTWKz6hKT/AJE+EIKCuEAf4KCNd5FYpf8
IQDGQvXWBTJhnOZlGn/JYPMtAnX1hd6iBHc1lp1mobq1JE9k0refImF7V/ziSg5aarHfI1kC1I/U
kQBouogm6sl4FaCjhJfcS+Xs5xYbiBKisVOjJSpBks21VAOLDmeH+wMp0XbKTzIdMJYx1D1S003i
9M4voS5CQPxXzubhKgadL1zc9jGCotUwskTzeIHX8vxFEyhAgfbvbHkKW0ISCGEC1wXy4O1B3BCn
zhEnvnFuNpNp1VrFq6b/76qed5w5MJUKkrRtXBeKroJAXydUmReiXuf5JBY/xRd7p2VSBF52mFqQ
dMHxvddBsXiyeDARjYvxSJ83T7tmo5Y9b0ryafwlRyifYRncrSk9Johmz6W+OnhNb/M71XqmDIJ2
o7bTauMycOc8Vq7vObAAUPNAJO7Juu26pmLk8uvXXGsC8cKl6GPgJLeTeY9fy9jt/3MbqUUMVDDg
bJxgnAOpbjH5z43rrke3gMGHtyR57c3JmBrAHyFPa3p/KN2zs6OoKK4Fu2IgbBiJCywrHtUMRcWn
OouZbe/npJBt9ehVx9QmxPsM5anHfbkMibUfboe4hP8Y3P+Nm6f8la1XDiz9MyCNPSQBY1AzFsLv
NUmfxKly8EEMjHATGeo1IGGqVf2w2PO0bmNyvisLsAvFc6rZTQRAciGYPg8P2WkGvyuXkiiSj5tU
VwBJBvUfaz9cvri9ze8nKrrHL8+B9Q8duZy+XbCp9TlGaTBSExxHsmo8Deb+mfGn5gUravcu7VHE
4dDR4XsornZ1THmyOZqme3rKBUKcFlUVdQeiwl4ItT23+CjZ35mXet7RAGWM/2EQV/VS5zTM2Ww5
/v2jiuWyiCZ7Fx3az68BS84GMP3joxxtgApH2Jk8XuobzLdNwQqx/wC2Hh+4s3vb7/LpzW1MKK9o
QZU2Oq5xuZZILduM/CW00kwi7mk7mSJdbE08xJTYCApfT3yzKANltgLcMN46SYzqJ10FDkJ0NQ5m
0KjH5v2PTLiMB3kYqfdceyFw9WI/NcX19IcLtWtOa1IskQKj65MME8S1QyAkBZyxyKSfheJucAuV
dh7E0g8XsXGHvZxXDWGn48vguKEDKBCgqL528FK98acVFN2tW2bpO8L+eNcJ2NVE6on9kjOSJstE
MO1wE7NOgTxIE7CSeKfLZ7gAE5xVVQVh4bK3DZy9jDsKKbapwqlpYj8sKs3avHL26hWmTq2MjtxE
7uh5XbhY694fzkWnf+YbBJJR/a/GqLhK0IYUTqtYM/XXFWppogp/NARP37hXUNYDqEY8RC3VSmsl
yD0rUZiAGuZ/3ZlX6J+IWz7yC9pv57ca78JDztq/ZFuLQqfAiHceCRcX9GPScaPwV1h/n+elEJKC
x/KUwd/jOVLJgBb3jwkiTsd7UeUnd/xFAM08VXT8pultAKG8ptxAv3gFIu4k1eofush2KpDoLr3D
BmE9b+pkShPygOkzZ53pFfMVDsxqEyy1mjgyNDs3H9FUyqGhSChvgfBb5aJbfXrpDvGm0uN3XjmV
ZVQ8wzm6EjGCQEeQ2IyQEzr/BDBOotp8Sq5rn/odFb0KJWPr+F2r2FfEsgME9V4BHnykQLwmCT//
ONJm6/8hpFxzJb35NZocK65gihzEu0qm+vn4yz4sad4cinkuu23zMXF1UwWZdNyp5KLFVdNH0w++
3BQv2jpcyeLW59Z0mETo3hc+mgOj7NYJtA43sky9N3HklybTc6pG3BrfxvtspEhxNjP+t2Okrn0P
Z25YUUQAwf1WaB5lpWZJyld3jGj0iA633qBTM/WyCUvbdta7qgpJQCdo0NqgUjHCgirw4h7c9hsr
En0ABtZuvFGJ0Sviaq5/cuVVdLbakkXLzyr+MvBDa9b3bP+d40D5/dszM3hTfohbsapOVfIQB2AT
1hoBxW5yyqMTFSZNgTo+3jcVNo95tnSvJrtSg+CIz1lI6Dhch7XurUQkngfqL3oYLmvZ9F2y8qpK
J+Df/MaaaebbJKSFOQDT8N/K+p6zdalE57geel/NHPjlcilmdwV3jxEqffoQevwJdo4tPVLfJPFW
mkymEXgngrxvMJjJbVWNOhF9FJ0/+Sf6Iv/l/fY+aSzGZcQiONzNUYLRwzAgipyIM7wl0okUHXMC
bM5Fx38vVULMLVFVii5ZgCMzCk33sVzHkbsha3rV3SNMedI5HPXJAoU4O7d1PnhvTfXj2Xo5KQVe
Uvv8DCPxVTatNt4iUIwVpVeiwISjewrKkePk7L3V8AbejkNdHq/JBW7RgNoyr63uHWZPpVSp4UnN
ouFHOEkazGcfBRBIkmDnKYU8yy0DBqaZmxBnE8TPiNQ0Rj7vV46QvZEORRo+WlBBHaU++So4Yxd/
dpAojmSL8z8BeSfOsxyyVA0nKVrZ9iSF4beO+xxvMIZcteD4GcuJQeOUovmRQH5sUd/AS5Gpe9Xe
1SPI/EPQJ817dS2gQtTFwvyvocEjxsmpG1FDD2YgDJahDZ9ZPliayNRK0mI1xITWQhpwcztBSX8h
xJCDzWMPY73YvVsrQGMgeK12FWgpJ7Ld43Ud0FrVI6jjK8wdKIVgtMBNN57tYS5UHLTCayg9somF
0CHQwIYdFbty2M1JpW80HhiCUHa+9xY5QnIs9jkvXus/VEKPgUokntOR/m5Tx89NjwqYCLTu+EMJ
djXxsgQSdpqb35HavujEgsGXXOpjV/EaQI0qQxFkAfABhmZeOXpL39FI/Pn2s3nUribWXbQIeAxU
jL/zpNhYGnZyFajqq3WVKUm1HCQEDR6uQscowJq7SNy1yMz7/OswgBMDNJMojxN5DGsOzUGdy2u0
vQWTRk/+TIfbhYPPPLrL4JE/KZRdvJfZy/mEq9BAjLyIC9+kJxOW7SYqEmyPfVKN1aAreEf5cteH
aN7HBQpbBD/mfPdMuZbNQQOiaF/gTQ+QuRimcorjgoKHZcGtj0l2wbKsQKMBC/u9SXJk1oGBX8dU
SU/N9mhoUDTqYsFeHj/G1WX1Z7Dsz0ZsB9LD8cxXDXIGBa0I9EQsajoOiwFpuVW9zDGCbxVtuwqF
3ExScb801fhR25apNiFVytehHfh/Xxrqs79Eph9dBEnlj/QCpVeAVA298X3VYIIGb2bjJ2pDSWVz
XsmZLjqy51qIPHQd4+azFuzcHQDcFxn5AmpaNpHw1FPDBMPp68gzqQv/wnUnZCBDUrZreEoIH/1w
hjrxgBFmtqIlPXyIhrET6bkuo+2BYodFZlvq4WYjQYDH1zKikOntgo8B5jXMPjpQQ0UdrfeO9XtR
oNTC4J60GQ1+IW9ZhyIDKr4vgMjSCrULvh2D9JTVdrJc5kpHgMT4iQ9uvjq5cEgT/Npfy1nqjlph
4CnS8oJgkHa6HzCRmlXK4qV6Q5QNTMA0FZfcIRvu2xrXA7YLvu3+SmnJu2ZELTYS9GMFUTb4GXVp
/t01VaSUcNXHcHgQbpvIYC/WMyoLk4i/HhvwYROSMNuKFN0T0w+bvUXOFPiyNITNW5voyRGRy4wy
u2saEtZT3ZNqHxidT3P8oR7NDprgg6Rhhrn6pumzHrjAUgsv1beD4BQNfJJ1dLADvlY5q8fSI0G+
8/rIjw2sN1fJOXm/rQ3NzE/aqNSP1Ez3fjkqI9Bd3CewS/pYqpDYrXX639B9K4Ecg2yjC+Q61cO3
JLE0VqZEtlJJLHYLv38T59LoxrVCYjqxpVNy+k3hMF+xjgwmpUB7CFd3/Tg07AEHtt7yNyQUhhLz
0QlimMFRH1YYmHXZBIFlYTD3DagbSZeNNQ9EXmIqaHByoHlhJ8W43B9Srf1mFUvtQF5sktZHmNHk
lF55yqo1vTKBdwdxr4RvC3mXQzbsepgAy/zl1QGHJ/wNTEdcTwDoeZIKFqcguUoNXqI2msGIwSsR
ldOIoKpBqtimL+qtsV3pkybpQ1WU+ujxjKEtUZoqnFfYSZw7y6+y4hJ86mUh23h4i1UgllhlIaqx
4IsM09QWKDkr6pdN6fmAH1/iKCFGTG2uj+bOzy5jA9INStjNlanJwk/xtcbdy4LDJzhDaSCnP8GY
9tG6M8dflkplPkkE9STvJlDzU+K+8D+wfDMy5w0CmGbMCOoCoI768Z4USaff4Y3rKj9viFBybKhd
l0Wd5GSMm8xioCXjjuFK4Z+XoYR9d+HRF9h/wReIR2rEDatsLfw6pAkCDMCDo43gggjUB8xoHwwf
N/dk7J6C3tV8etsXgg4LVh4GIuh1xbHlRG6fctDzKm1gq78VmBU/oFmnw6Pq7VURyr2s1IRI0SaQ
C4NSnGAX58SsKKU5I1mCPPRVriBxNWVLn7+/3sK2cYjKWZqBMjQU4dVTEhUIzhAP2tzLCO96fdhD
XAWBIEoenHHuZcJCpt5oI4sLNr9s5YL0qpqSkVfw4ZLFhkTXcThFCL5pgLx3IBXIL7BVq++hUvo8
h9+wdFYDenOKlQvK1P3RkMQT22LpLf7avHUYNv2etJLjfb6K3sx3NoanYyGElcCsWfOasvcg16eW
/Y1Q3GKJxuP6OalBq5FZ/CmtOilivz7n7y6lYeIq2WVmBhXuS1oQIdaSZP2DVmTeTEmcY36KbHZg
ZNTt5CqGKXZCJQTKluESLSwfQ4xEXvemS0P6O/mL0qH3pL8NYTnwg+6H218nqy8c8/YUXrkS28Bf
31dQvX49r/NDpTo6Cjqf6+6hvogKxSm7DvAzNmDWV8Ttuqfw+yG4l9vI44wnxRcok8JtG+ceRqci
mvhckxXehMCx6shT/rIz6a5ue6kL3S9nqK2+lmXLUmSRJiE0Eh5YmqcRxvowh6FNbaYBPUr68TTr
ozk0PhvmTMFyugKwAFHhcImbH5wIDbOAnc5oIGeuu1C9b3qYIroyxpD502zkNg20YTAufRFYQbcw
SYq5cFf/c0SqqJE84CA/PmpTCphILb0SfvMHnDbSCsNqknjKiJousfGvDAvAJbbx1QYG591/DZE6
kffcoN6AAE/5+VvqB1jzyOFl6/yjXI6hiSInC5x6PEwuugvq3pDw+MF/mNc4ZiUEpaHFd7ZMqUAH
v/rlqw8AsccV2WqHT4RvytLmXEsrwEq+P9qKn/lf4Dr0RGqQzdWFdi/5rRl+aR3loirwoweME2vX
DhYSTc3A44T8PzsrFxHD6Dkt4NTwMa5VOzoGeiSIpCV5K88QcR/xr4Cpo4MziwmhkcKTzn2GAs7Y
/2sZbNKAPDZ5VShNflhPOJ7ZGv5az9UBOUs9yAHOP30FOUQ8Q2uNbQTmRx3x2AsVT9tZrGxmEI+a
of94dRM+E83OAilGqWvLY20K23XNgW9s963YCf3j5E/Jl+iBe7EbkkoQf0GmPxW2TcdhyYt/nAyO
zcSvp4+Ah1EOHo8Bql8phM1GQ5LKN0F9u+fw7FI4U/zwpT7Yk1qbBDEuNHNVC1TmnFcKLYyDxhwt
dcpCpcvo4EL7kk8ZzdJr9fR/CBgPIf+QU1euLEQyhkkdxFgzvj9kpSbdpTAwmpfbbdF+/lJFBiOF
TiMH9A9BKSJYXR0SlmF5oABqbfKQx48y2raeECbdoBxEwsJMU71Ku6rNC5qY4Wfz/zaNM379qEY4
WcOppqa48vFut/b36BS2Bdyv4pIVsUBOrdk5rM1M3L9tJhhAndqqjyB+PheisNkK9PNQGEJ5Ylwf
6TBG8zgQalC0Gjwgx7eHRACBlK0F4QA3DBlBLosGRX0hrJhgfbT7zWV4aYXE+Wl0Ly8gvnWzqbNQ
lw1aQ6OtL8TrKom5bNAX9KiBjjpx1SAkdyPCEOxqPpViEswJNxUIeGg/f2PqoRBA/ArYpLO/A0AS
IIZO1jhHlSkVpM7MkWdsaM9UKfEDgI8MZERwm2jEmRsxcRB4LM2XhdKmfQElBvuxUJqD3uL8jHbf
9yQfegqyaTgesLiBC6rg2EYgDv+JPMJ/bsrEDSJUXOq2pVijn9TkLf1xmiibxmDKNK1NMMOAFAuY
d8hWkV1dLHUcsylJZkOsUDhV6/l2ZcPoTRkE7IxIhnW9743NQmxlG1CW5tDX1xitURWUkGkI+Zz+
LhnaQou/NrNvCMMDsp4YMhtl7FU+HdHbgnY8lMm60C6MiOSxMrtKtFl6gSZs3rFmWzZeKj2qVUCW
mI+uJmr0bROoPWGUjzdD14Lm5SJzhnAxlJM2+DiMCjVc+LmdCZuv4Cmyu+UVGjfK/xhYGwuoiKmp
juqWF6LBoLsUSvYGjxG/ophgfVbt/sotd/+DnFs+9ZNgYRy8W9A1/XxMVyjWkGCBYqMgcVqkpNqY
cDYPUcrMnHLbQPvqh4RzmUIm4vAs9DUocBDSA3SnY6tYVYZ5jl0CLFhWtJoJtvv2DQcbsTmrY2Kq
z/NKoohcMyNyR6DuHDoCp6CRHKHRNQJkXDyqh1zPpgPXJkfbtiZoUw/V04OtsTLLsuqoaWjCDtLv
5blE/DX277taGv1ndhcxfEERnbCD4mD3oV2eIXmc+LDE48IYxBBDH0zOyHLzLteLoIkoEsUVCAFi
dlAcv8b73LK7NEZD7UE8KAJ1pU0kSUU7+FxrUhm3KXZyJDVfAClIfBV67uGly86Jz2+dOEo4X0QO
xvO3fQU4JKDABYHj0u7SgD2BCqyI6bRfKjKdT/q8d7Q/YgjPq+eA6B71XojoWB6lRUOioE5s56CA
oCdM9jcn8bMmsQ98/H7oC5wjJOduZZVLlTikDkAAoGelN3BlN79w1tElfDWv0jGIgGxOERGBBTWL
zPqwunWhG98UCRSIBmjG0k5P6ZzjdNYV0uVabEd01iNj/qSkzlcfqJHATc4xrxBaAVO/aLCrQzrw
AQd+Y3yyt9QS+/I49wlPZwr0x6IL+VEzjGg9dWcoAs31xyY9Wd3V4SFgNBK+cZbQIQzkOnMkoBkV
eVMLC0CmcSfX12usFbyh95L4Zks3Rv3T5ZlbBp8q5R0xJVDLezrwIiVRMDB1Yg58sFJaGsmhl2+L
zuFimzQRcW/AdV//x2gaIxORUTDMMD0851DZrRyRWjSkMkN+VV2GrzyeKGmBI1ubcqd7btFP88N9
W0kg/N76PHv0I8WXXuiZLU8qcue0cFb+1+ZF1+CtAjBFXkzDIlpE4uZ1nHpS+zNY4MszqpXnv/s9
io+EQ7amRATjT/jccCnt8IaCtw059wF4BJrVgas5Q4+063ctTsbyv0mdIzDR3FZ828wy80j4241w
Lee1FymSwCmFr9LmzkCgx/4vGql+WwPmxct+Q86PbaZ/LkRyv+QvBCaAvxNJnkIEo1vAAv71qtJO
wUeIvCfOBMsogAgj3gpaV/kqgy2don9gY/aNHDpDUpnLy775C7lNMuQTum6ox1mDJu/WtFYdGZ4Q
N4qnggHVIw+aunRz+SJkzpBrGhgyNK68sWqXeZwFfbgH4CqtU45aUkg6UwPpmDqwk4FEXLgqrysC
pODkVM+UVBwkqfBSRfLp4W2/vOB5FY5mKBHrjGBNqT1WPCUfY2RbYfvceTq6xmKtN+Guc/Avndo8
sgcBMJBA2BDA5Y9EdCa4LNcqowGvlMzEOtTorSS9hlaNNJtBcKvWDmDJjOTpnd9N4EWZiNLIeTM8
agv6aNLGz0vJxzdFCO/gtpJ9IGgsx6rN2vzGBb4IbAHzZibW1YXcD27AjIOHRLheYGvb7Y7KrEkG
2i+F0DSFrV81aW23A6aViqMfKOkmZBjStECnVK8rSRNgxxoDO88LoCZZvr9nuH7adYh4AVA6C0mQ
8BzB0WGXlwZsp5bIXd5FgB/AH/ZKMbogfRQDvj9vxxQmEAJC1aS5mn3NnIjD3r6MMV01gJ1Gaokv
6Vx1R36WHZJZ+ceJKFfWTHcAxsqYZrPGo5vz2s7J11DL0NVYPDuBke/wab46taXQ7iZKcIZpHYzw
4AHwYD5O8dofGNaAtFi54J0+DlxzZbBl94QJmWAQZGkjYVL4xy8u0htpGmbmRM2eaOCMpYztf/dw
QXS/mI6omJbNukIIYvtDm6Q46Ty+kSWZ7LquoUeTcT88kAOiUAjB4+TdfVD80dQcvBMSZ9m1Wgcf
po4PrQshWeBhktjXBv4+2cwO+B8l8AEhmkeB9JeBdJI97wZKSFcF+f463SuhWtySP8kVQSHaGQ8Q
ocys+B+vXB87LLSc8BZH2TLCMiU8up9C5mKGNs+UqmhY89nObO/tmAFXxM4TKMuomV3Vu6lSUeIs
UN+TN9Fi9m8S4moB4ocfWyLTfZBCXvNWQD8KoozjYq8z5htcFisf+w0EuI+p9at6f+uSMeqjOvyh
HWV2qkdK5geESSZ9h15kbmea5WCk+A0VHCcMIJLsLnkWSUz83t3f0hRFcpTOzNny+i3d1S1re+EP
r5oUJzlITCuV8sDKPrZJanbozuQecHQLmIvK2p1ZHgorN8Y53RYpebK47qYI4jGK8JKj0urFDERY
Jgbdsa5qeHMzNJq2t6HzUZ7gcbKkCII6zE93a0eqnUkte1+OBK2qIDHxZM3evinqZgmnFLILB8Cy
ppctWXCpCwB6PDgAM3qG2OWeSt0YeR+610+WH1ntQaKJEdauL9ZUSMU3t+usrNl/jt+Cbbtu/LTK
oT2rVle4FIr2CEURIWIg2w0Wtdo5izgoI6jvX7MImLRVEvybXl4qho3NgZegwTH45QB6QTOURja8
R90mGm41Qm+7pt5jQWY74aB4oS6OngtLjaxSUc3a9U2tsPnInpuW7xHoOGp0DntzNcC2d0OOo17W
X+tWPYJ5GwlrNQldIQToTUNDIENaDQe02X8IoUXJYYFvvnnygGbwjrmYXDE2Xy6OiL65xjZ3q1yV
lGe2hrR+xIwUsfDv6N/D8iYwDoppJrCX6jSvVETm9k9CuV/JIM8v8Pl63Ks/EkwxirSjWrUoOOOz
leVRCtkJsn1apaBgpqb+rb3j1Ja90FmH2hvqxL0YELluZtbjcSxPR1a0BscKLjZY7oKfyfa7QmM2
bOhFTtvNsMY2PbUEHVVsLxCKoPmX4154tXQSc+0hPQiIpnQ7H16WjIba7qRLz7pUDu119Si+1ePF
JNA+PPfKE8YaqPsui1toxydv16dw+fMFdN0fIDTVpL218thx6EBRTnEK/dbhKfmy4LxcDg7jcbQ9
ufh6umvvnf084UwYJEp+bpnTx7x7MQtUGshmEQxdSxw2NjbWSPHLZbf0wmC3ZrGCSSgeTAZJUUIp
nMr+wv0z49JQ0fDiYXsx7tOiFyOqLxcnKDaBqFL0EgwT95UQXevrcF4GWg6iwDlcru+wuu6bF/kg
fcHaXPXgi0/x0apaW2EkJfTkxINOtlXvtzYlbsvt69nUt9+PORd1taDh7/haAErtSHfIZkP3NPtT
OVeiwdleKEiZEkhDVw0feDd6oBNkMy5gXlsGgoP+V7w0EzhtSgGde8B8LrD0ppP61XG+QGWAK8lI
P1fUmZ6DXQLY8Y2y/X7OKVSLgHdGylmqOUaTjV6CG0pWagrnKi+nk2HnZFD5u/PQghbMUlb1VcCI
BIyFOdSJYhd5zY0uR6MaEpvfqwiPcdSnmA/JjYuuNHa0ziZAE9ChczlSNj9fbMuPSl8dkdtaKKT8
vY3WRgnjq3HHvELMlnieQ8lSvH96tDCxB1LcqfTlhHEM4YlLq+5PB03ZtJH3xp7tYjkvAi8/F5Fg
LGXF2Mha2F+MxNT2r3Fbctv1J2Cw45h83kizkJODbcug29RHVrzf2OGYn5X8arD/xtMIyJ9xJaog
dtiONErJYU0sqX0aCoPGruW2Ltjd552z4TtycEwMkQerovNQg1wR31RKanF5QB6hld6VxuMRU9pN
zaTRRIJbg+WuWvIRa1CLQ8fLbiJLOStxaIuquo39MP8c7v4VxNlfG9QISLESxJx21FJkHA2G5ah1
QVD4g3TiXl+ZIDBhkbfQgdmvK8jFZBKv2yG5PRgqH4ZV62LtzEZ4danfcJFSg73N5Z8M6EMHMmN+
CbFTvfybFA65tVjQQxDg8NxUwZeMcTRG1sFEcrP6r8XEMSc+C9yRZvogMii2Br+jXS0QIyIh2xvq
v1x/4LBggTcQp7vKhw5HbkVcdhSRsNjnHt9391r0wlW3x6mhHnCJkt2CbE8YTlcc7cgKPSvbxr0m
ISTq8avDDChEDjNWyE5w0tDAtkKPDRs/72YloVHquQbDKZrnpwmucXpe8rgtsTFQaaYPvO9En/ga
mgA/bmBNb7d0nebPvPKSd14a4B6pHo7MvKDAXDieiYNa1c3KvaFTDx8GY2QX/YhwYuxQSSReIdX1
ytH2EiYuxhn1qQI5Ts6MfSf9vB1EuFztQ9GXdCvvzk/ICaz1LyA9YG6PXAnkDYX31Vd8wJ7ITJ3M
4P70vXcCEEkRpgWhqZCjZDyS5hSBpVHZEMyfdRRd7oQFvXuBOB4/+l6rSgNhrdLd+JPHVgCuSGJS
ZGXZVaiZORYzzf3bBnMK57skw+qt36iqW5yhRvT+aV5keZ2pCmVMkjruH9lQbaBJ9WEJgOH5jkXG
6akEQ0YSLQIeXB8rFZSMoGkAE7Ra7pVyzBIy4cS+Uzbosw/fEGH2NX/OYAIx6U0ArxIb/64LEIoP
pu2Hs7+u/KYnf/ip5GWPt0SgO9i9Zz7Zpm/VbimrFPXFuw5hr+uO3fXAEFt/Se7P2CPYei5GVc5O
ZVgZuhyqkZYS7Ojz1jEV7qemlMBEE2+regf7PtP50uu8zP6C5AM2dZtHsGgQMuFjPlFNwWlO0ltz
bW324F+vjOyP5GDQUY/pfon6z6+m+ON3rS7R0I1pf5NZ1Nj/GHayyQVeyG70/95RGq2MtAGkqws4
tor19ZAJBGA8+t8kzNFI1CfaywQBTRcLeWLiTxLPg0rrhU1JFrexn8YBttQ/J1PzWT0J2sVvKwGm
78DxTM/rHYjqUjXRkRqNjfkGBlHYwQIUXkQxFUx/vmJJ4B4HmwIpDudCM3d1PKTOl6i6G3cN98qi
pBHDm3pS8kmYW4aqwcrUWaINVFGxX18PTd/czm86HLsB4/wU1t3refu6jG8W+mdmM89N6aFa4fFP
ZY/9T3jDHIgja+k2p6+rejJGgHv7uCDBqlPx9dXrc91gjHhA67vAQsXEtda6Q3dSkfinv9YdqVb2
Fec4A7naIaDTUg+tULyje7s7eeJoRCUtfrFQkBIYlMKwoM6GybwwB8Fqk1QIAnKzBhXoq5fjRZtA
w5wIjyxbqg5DwcoWgaEbeOWvT+rkHSKZmUK08PxL5JJxZ4efBG8jfEZkp72bjjgqrE8pppcpXABx
0MxLXjo2XPrOrxp3DcD7aLGokv9msgdgTcT4GLU3QZk+ktXKjA/9mL7j9fK2NAA3Dh4XGat0vI/O
yrLBe2goHm7Vr4CKZhAvQ5piU4i+Zl+LWOT3ZSe/PMs1KWpsu5dnfTZWU9hVHDn4X14/g5jhJxb4
4bOYguoCRUg+TPS8y6kHykA+qxIwHELrsiaJzlK+FJHxyzizvITjeBMBNt9DAF6lynOg3g1VZ1w4
dShKXvandHFG/nqSuhXLwJT4TE+qDXZydNZtKRt0tbk/kqdkgHzZaEEckhtgpqOYmCXvTcgfCU/q
M+oGZ+E+aTigy5D64gMEuv9yP240V9cOKyEA6Inj4VEl47khoklHK1VbESjNgPn1ByeXFcM6mjum
ohTkLpocdUdk8dvzMKH8HCimZXv+1NSSGsOBAx/yazW1WiCabxnJWib34SbKj3YfgN5CHaEW3hVy
fL3LM6DhtTdscxQmFHaRkWER2s3KEqFZrACr/tasqJp5s+hlFyoYfoIpYoJ8IBd/xvd6BEAi4Trs
87cFnXG3eQT9u33Pb3XbyLXrwiMMraxgc+zI/LShmxsKWFg57nR7Mou2XavQI1u1r7Id8bVto7rg
eyXRyHvt1DIchVeXvAVLXlg+gNxiIpaaDfjS8tME+qdWOPrVmeCVfgJt+s8PmVPbvbxzI+yljtpE
k+U/jp3d0f8BY+Npg5TMzKUHg3RYIQsKpIEfqwi8vQnyQxTe1WU1wc0fV3iHCGHkj0QZVaSbKMsi
MbRIVEaObDTw3jTiscEWEhDk9AmcuqEjMnlDR+p7tng/1EZmQPiQSOdOdFfSlqcX++K10BGHaI9f
vnsOqLZtWxBduEtquWzwvDh7z+mbTpWRBkEuReKxvy/z/3RTJ3QGxU6Gjn87HwJz1F7wOI2vUC1i
D5Q8kIY3AE+3SY2X1TzYt3l9kQnBFPmeEwBlTpnpuUKSaqaJUVVTXu+hY2LXnGHgiIEDq4GP8wMG
0w5hcUZecsx41WJGDCSud6FWHRyXedxph9zfi7ausIQUYkG1/vu5GZjIM1LQhfQaT9ZT6XIilTJM
yD9JJ2jFVNERL7qA/XbjlIfPibWqpc14kJs+OK9dMCsAnArEhtusHzzJK7Cswpzr5xVZ4NSz14qX
AkCmnRo+9hnRPDcBDSI9/a6q+0sENbSRsMF95LHw6Q2/Ywynq9U9Icc4b8pkTgGvHqcRYly06x35
mGk3Bs0U1CAnDLUJcJSWx4A5PnD0Qi028X7FxRZ45xH4vKWn3UsoldkJb+sncoAjFHI9YtcA2DRQ
ObpZPvRQL/GhgcokRm5tLWhDNTlaTM6cVQlLocdO8kEF98zxivb3PBk0Aln/fdptTOfeFKpAOvCb
H0CwHr8XRwrjBGWT9pVzFUcy/iV3JJKKMI7MNWg0G/Wl5mG4CO6c/yui8pYkyjSVP8CcCSS3RlYI
yuJDxiIRzXJB1yBZC5Qjrgz/+rzugjWCIUGPJh3AV1g2t6j8ZPlC2cTfJ97YHEP6wA1rQqEq+4O5
IBK0i/L0OuUoCLdRT+a/J/sdUzxb/R9ZoVRyVjo6n4kcpsVBjhaavzAfm/+IyixH+ZO0n1nbuZDR
eaFZay4bWUb1hwy1TFvRvqzFMoFlpff2HfmIyVkiQKhxKX6m5i2KY4va41trXmqjrsa/BHCUaHTH
fmn5rTr27ib2EI/DUFcz9fPT7s9SIzW//mObdbrs+WWNEM6oHGQUJV/Qh/KNstxZmZ0kdSmiECgR
oG73jTlIhlmkBjSAzCZ0jPnup3dOm/as2I0ODbAZY+mfMy+U8l9W1IiROggIzcjTRsBsFf/GZu+e
pg7lgOCiNYWNciKIxOurz45NzSz41I/i3jCt7CIMMhoTeuxVE1K5/Ux5d3wKYRzBQPXpNQJv+3yv
YOhXD8L+JkS8vQLFBxvE6P/7v53QSE3NZjmb6/MrDDlaU8hA+nbfvNqpTF7HmHkosQfcQbEp3A8G
TiAtmFEtarI+JvvhXeUzakAVVNXL/ncLLC0sita2Qw1NNHpIAUFEePEqUA9lQTgllEIN78bUXwSM
JMUYNDfR2fSrq2CKUR6M1W9TqMngC3chKXoa1QgNUZwhqRGehv9USByaU/LqVIlTfhM7UQRcK6Yw
iT5RgLvvrjGo/iNdIwkuc1ReUNuXvpGxUGalOFhkxqXQJx/yInG/U+C0C7PMN4vXaDqSPHtrZzAi
4kuxNEBfmqVpD42ncIEFhgXzB/rvp1NbMnUZQWEYrDVQgNZ+NgvDtb6cW9jyFaWyX9nrY0k47R2a
Jm4XnyezrYwuo+vJvkjo1Wh/k2Oi/BurXgxpkdbVCRE7LsrhXvYzSUv/bCRjdI7g34DZun6TZiZI
zhZ+NokzJhk+4U1q6dRU90pLkX6R7y7ST83tcWlUrE0goPTRsmMxXD7zAVGUUSjiO77gbsVLfIUR
BS5Jd/b4aHd42EfnYONPxuyww91D57dp5Otwv2Fz+PJh9aNPMShzwbjaghxl0rEV6dco35PDUvtF
mt2TkmayyQb8HmSHiLgZcCZF/6MWHdICCsMgowEfk6ig2rRItuhyg0a5ayTd55QQ0s1whFvXQYtT
Ot3v4rnedGKUSzo9GZPmDH3uIfC9H4tpGs1uLVJp5X82H2sQPPengkz6tB7pfgK/BltaYHaMSYk+
R+l73BiXs4Vu3AxTeaV1kwRKClkeP1qnZVnQ3WeY+tUbx5e40gw6DivAWWHLS7vsc8HK4LOdlJu3
GE8Koqqd30Anp8Zeie7gqC2TJzftD04McbwIvBKV/ZRoLearon6DLSc5E37QFXIbAsQYGLMyKiKX
jCTxW2j3diaXmNZyiS10gu/NZ/mt9UgqEWQvi3BaeWYL+m1gvew461zPVKfgUug9KMqjVOUhl2ma
GOJj6d0lR7K+0RVkwkjrHo8+qQGUHDnFxlMCJq5WE/+587Z4DvnbmT6NpIGUs5EQh9X1Ey85Hutn
4Dbkd0KJos2/tzW0hw6pVh5XkDc5B/hP1EAlVTD8aZVYpJfW8Q2tI6a9JVXgh2iN1bUf80BuCo5c
23zaBRzOaa/P/ODszwXwYOrQqEZ9hXIyw45jbCd0qcu8L4vyECQ4D2nVnz6XUqklZR096XD/iuHr
/z9Xv3dLBImkiGLmUCV2/9wqI9Nzffrr8d8kYyL9ohzRLLqiheLzoKFQ7FM2fZ9Cs0oWgcApllBs
yges5y7PJvr+DjPnCmKDfP5KSPCHBsOF9sNW+GAKtf95BpExGAz9Z+Q4d4by5xcWZtmfMIqAd3Y3
AKKIHr8m6KeYGF+aMFwzgox4RakL3ARb3jhipcwjvyT/WmVyAcvkkLFKmhgL6q5ypuijZU1KDobx
MSYScTuOvAoBmUtYtTLOjuBJqoIruCOKa3hTDYkXJfIPDv9+gUq8DEBrXI26+K9/sJP5Eb+aqQA1
vjNTJNTnyBJ5ANOV/i1wSrTPhLbgTadGtEjKSEkwm4nOscAeCEbh4JajxO6U2gZq5BrSjJlIbMXS
Ogyf5znXnwloN5EX53T7jc8U4fK8r/DDp5WJVRkPGb9gsveFQuu+FwXR11kL6S0hk3YZ9pSOa7Nt
zTQe3+wC3/LhnepjfcyIkIo9OwXYqhVxzmk1CY4dTQ1wksIfPIx/0HFFEiD2zL6uCtDHFun8bpxZ
Hur6TuHE3TXh3QC2swCDN/G0Jet6WS3+GbjsQkY70qUSRxZuDHGykLZyxLC0EUXKAXKPOmtEqAHd
KhwGmbDGoSh+7/NkNrcsRE9rANzkFLfVDkQHn8jJUeO5SMVcGwBRgxMc+S9fPch/hG1EfRgsasMY
41g3YlZyOkb8nmKJ9OhGgLgFQn2DxpKxIkFG+I2xx18lpSw5Xu7nFu2al0UquJ0xZzarCYCwezBi
IPoju/FCg0luxP+hzAPiFubBRv0Q330Y7+IUtkfSZJLxPxtQZGj7VgzPSGzUjtGEuoiUqI//20f+
Du69Q/Tjt/wuqHFkv1Rll9icXThIC88ZRQ6r13yj47/ZJhI4Lm3PiDYDYaddzc/S42mHEsmt4EQJ
5+GCIFVuBsIMd+PKcUHzOiamOXuB9pMRJyxmDPiQGps3PFqDBZwCjk5BFf33GW7l7Kl07zLMY+B9
POypjzpGOMwK2kL/0B5AqPcYt4O+lW2Q33+SOaaLzf8tH+tTTwElhPo38xxayRxPbgbzyOBCZHvf
EAgF5NIJj/9pjsbt8s75cbUuJNvLg33ExA8qC5srv8jy/pj/1CiiWNJLZYwYbGVINFa1IcplnJcz
ufjpA7nour8HWi0U5UsgQEI+hm1roO9Nc+KtkF4sksBPyLLx36GwBugD5NVyBrdR+Skf9QdqdgqZ
+AtUC/n3S5F9VeD0n9I8BB1k8SCeb/3hU5gN272BUkcvD4tBov0qnJql7zGH8OGzTMt/Ol+bK3Kd
SK7LRJZ4qOXNj5j5A8moTT4xJh4iDLrPVJz4g9NQ/Zhbo1FSkScB6fcJUG1YzHWlO+ej6HJ5qkEK
qVfk3BVXr+4ZtJdOt51M2y+4cNcMs06acQZL1Zf0j2Tho2kMe8ZdwVGj+kLT3/9rtgh0zH1z/qQ4
RqfmoW0FhPmZRPeTJ1mr9yVKlS+gB267D4AUj6XthW/cTlQ198uzeYW7Zbqp+Bwc4u6Gvzoci3ld
1Z9LEqgSpwXNv9hKgRqtUONRT0YTqkQNKaKnk+s/wIqKWPFOlFbhbyYj+i7AQOrJ4bavRJVDZlMQ
t8EL7br/sJd0I5R5aaMTn/lfc31+TPJt+uaWN9dcAqXo6bBXR0+fbvknQITuH24OzMVzhR8jXcUo
D1cV8Kf51E7YoqtywwL/4rNH1lvMFozXQnXq++mBMp+tMZQ+ins9W2DWkNtNnRxXJ06JtlDXwyfM
pxW4ir2hKYGstZxdnbED49ytggvl/lEgSBvZe8CBVmuK2AxojxIAeBSjb+f3Po8EN4GhGaIWQew/
gKr8kNHHzfbrgod64PkqSKFStNbj3aOJ1ODf4vc0WsTn2oW/K3bUy51RPsINUQqwWyLMQFtHWxsd
O1nZSNlYHBgQjfH+VuIWVCgPu1ky7kVK/Qm9Co1e5Y8xotTVxfa3icU79bg03IJrRg73CHQncCB1
REe6gJyKEJEpPOZ5fyF0APBgnIP/obqkSIE1eEugB8AkLuaBnJrwr0FtP42qikjVmKCCfTziHr2D
RBcgEKjv7E7frRrq9nAj9VPidOV3G67p/EGyYhRMw5Q+ZOt4DWHBg/XklY2rOtJTMG6KYEGQoy5q
XpoEOQlRqpSTWd+FDu6NCWZxrAyPuJ+zpq4FQURLp6ahUfrZcMREHPNy9b0HHwnUQ8kRjaQ0AbzE
btxmd0emx4WGrwgotKFdoOoiuwBc6IGk1B40lXQ2SjeSgc3p0E6Jgtr9gvJTlIBSLOdzr4aBI5X6
Z+QBfC7pDeyqOYZStl/Pvz6EXb+DEFccn2WJ3lxw6pGjIRyyu+ecjMkW9NeMyhQpbvKW2Y7vDSiK
mlLZcnNT2zHAoJcOHgFhaJueXJslmOlA7FLWc43nmPUzpodNXY5L2Y0xsd39DEiZhLaZbz/GyamG
ocTQ/xCc+u5upg0ptreIjxx8TfiAT42L9uYXYV1XOTq+9lNmR3hw4QXNlVCd/cIo8OAws2dRl5qa
y/CB4F/0W/lHg47cwfpyu2rUmoihdMfdMUz8vS2jh3i7d2m3F0cbqX9Fe9raszdWBrDLFBTZ4UAi
aWv316O78032Z14ImwnrIqisZ2vvVCisYbEtE9+1LBZL9F7wu691DrQIobbBfN0KR6DNneCgSFse
Xe/bWsYKoZ0jT95zN8MeN5IOygFy+bE/iBrodqxD7FwtRL6sTZqtIPvS13m7eMhz7f1KciqVwqv0
pvQoYdJ/+7WczbvGTz2TIIdZBF1pNALLElnG3BdcOgYE+HMESVxyIENpd+QlppALBy811fcgdNPs
LoIWPzNgkcuq8SHZHy1QzSGWOLJa19+PujmyrBZpsJBE6/lyOe2FK1ZNKG4TcFv4iwIgav1GYVlX
v24mtcA7+WYL+HV1fztlXJ/ma0DfL0jN0WJXnSBhExCd3hke5S9yJYc3RyOHQkPhOGa0BHDVowJk
ly1Mg5Foi7l8HfVSnBvfNrvbP01Nwu8i1GxriEbqOw7420+yFM4dhEOnklunWEL6+CD4G6HmpzPH
v0cu3Lnqjy70XN6ZapSdvEXqIeFEuorKh2rnABLeGznlzvnGhqQN0ABrt53nYUV6OKmwxyRUara6
Bk7KklBpZr19+Fog0I1pl6F2OpAnCp/P35T1/xnyTW0CCDDtQXlJb4CiC3LriHSZrPfjIzAvpJb9
8q8k3II+jLlGXXGCsm7yJGq3XhsuqeKRrVv4jmoZUmpztiHON2fQAIra3pQyR2mTaPCMdWIygYuo
PcUgd18kmlzhiJSVIF5yIW2m/FqCp7mhL1VSmPaQ4kNuLX+3H7amrF3ABrXIzpyR7gmDKWlaG9Kr
7Tj3AxyD8ZDr1dVy/p6KOrbko6/pMbPJoz1vAdcrLRH8v8Mzz1NguGAoiSo0f+7iNWXwGfQg458e
OGzoosKXAjjPliuRg01kkVY1kqIo6zltRWM8LkBbVOvL4SdXyvQ9ldO597SdgffpFzJdjKmq38kJ
PVByvIeKG9fjLLNMSa5ex1RC218fKIZwXA2ScS24eBPvpPDStp7G6bvxUI3QVmRQ56YJRT1q0aVP
dJAGwphDuAlWSK3DnhEZGvOyre2BMOTxKMobdxeHZrbz9h9urUA+PQOiv/al7iPlPkGR/tkFj93S
6gpGTQHVPu2GceRLUuvDaVC9cAsAOQAjwZGXiZyRKQlNPNfbAusr/azGEhFcDE56HRLX9TIA/rXs
enj/49wapLkNjpYZuL6NBoPQ37CApTi+yud4XrV+Fj/ibyizCER3JVRyRHBKw11/R1iY9XBSWLRK
iYO8/WVh81DK2ZAIfJf1SO/tKkAUMgmc6Aed8rYmwx0nmV8J8wkHaTkoZN2NWBgyQhDyIa9lVVSX
6KjIGD1FU6nSsWYGtyrUwXETWaDHZQGq7Dj1eCgciP138YAHkIS7s0N7VbdwJsn03BOuaPm3TtvW
1xqmhp3bJizXpkb70uEQfxU4PSAvzw8y87H9xZJCV7Syy6eHXoRCQUvj10iONQhNfWH5iYxYiMI6
9Htlt77PGFxLYEgkIwgQ9/eNJooaV+MBdG8CPg8U2D8aEwMGXtmT/gbPRyfyrWwG1Gnn4iYAiEJH
luB7EfA3m22kfVI3j/Zm+Xm9Rdh19qgXEVIYlu8FgdrvzCZ+wJvTtxp3Ncwpuil49DtT88QPhLs8
e44gUm1ZvXTnugAYL0DqhI57k7UFDtwo9GTAkN5zpp2seh4S0KizYP+xHSboGF0MAKDe4se4i2NX
5y1OcV1/oehRxkznRzkk6JpT2VCNqA8I6iPW/H/t7RAPeufaF2hutlKLEdDQTyvCGBac+hLqyera
0P6i7UEL09iWMP68PeN2Uwj3sVYlsk6PXNYBqIAJtRzv1BQs1+GgvaWNrW7nHA2MVs9KT5qwgA61
LSNmPUIk9FWdKQz9m2HBXzEywkq7EZqyDbwLbwS4xazBbZGQfBpU111mBuYzOQp/ijuGd2AGDWLm
5giP+/xpvFFKL+to2AFPwXI8MttEwgL4koo9sxBpA+tPl+qAft1w4pBBBVGRlkctBw3lrdHsTAQw
nlo4RCliQ1yT1nIppSzgUq4TpVL5GGxMoififm5Ps4+vQw/UonawMSjJ3wUf64Z7BeWn61jBwaGD
lSB9D6ww8/+aiCkR9L4VIPwLb8u0dZqwG4X6QlDlzsQfo2y3oF3PqoeN1gIMvLzyPk8tsxSTwKrX
l8Xiti+J5sjT9RG6vuJ4YqTwZHzde0MGf1vh5QFPFRR1R6rb5XXOy19NnVM8fi7CgsJD24Yx91TL
KIpWp1Oqi1cZ8j1LyCVN1ymerZcaiJyqKOMi4FJYxNkNGg/IjhBDu/+/Hq3t8nSStOfH2YSqBEdu
o2MS/OnS/Y9t4Qvy92g47hXRHKVUxrz/Ztscy6v2p9g+1Wd5NiGr6bye81sNYjhEZnNlb/Kb9tXZ
tppFqYQgQ136+TW1+gGwyNjtbNpaub63tKOEuKmV5ZI/NPj+16GUl3O7b8zFu+op/SvpK1G0uU91
YbUhSAwYDGFER9I+WzlRTvzGHT4nD/RPsoOh0hXgONhW5osXOyqaWj169X0O1GCdK4H5bSZo50QX
kR+enoICM4z1ISgTB7GLON2e7StYWuo/tFYecJLyFiEl24Mgb0fgb8ZwM1o1LY0/TyFQeOxu4u8X
YKPZN8sUDqyF5d1PR4r8tHpYSs3pvT+guZw9PUs9m3yFXcOHozx+bLyr4cMSCIBgt0GyuoW6bY1n
cB3ECiNGUOE/7M6ws9IH0tZOs22myGNtQPqyahNPpRq7PuzuAmDO085rXZwKYjHh1RodZK1zNC2G
51lgDrrwsHqQLEbVMoQRX/WWfh+cVH2bf2mMasyjGNqf5numkh1dU5AOXBMdaDqSkaHyNKEaSvbE
tHGiK7RPvgw1E2Kiye+YawhJDTcL+wT5QTkqeaJw8iU5LjQAMQffRKcpN46WtKQNm31IFlZSLn8i
ZdyBFtZvc7RPO0qgs03PM0tUZgueLj5U4YjDQSeIqNw6AdZcLuRn5h6IUfxUKrlb8fWkeFn/iXDw
KLK5IGcVRK+KRmqwNWOLVUpO0jV/DKbmp1DshsLSlnvS9EHVqQLOKo5O/PE6/0K2FmdYTYHTORbp
AJt6xBPXvdtPCnG3wWunj7Ahja/VgPD+/wsz7TT0Zk62ZSNAWXFJ4egghmzXskI6BfpyjNFGIXBI
N50mrc0fpHHeSaP1k1D0vSOk/BaECXlWaDsqQHnwUXrdv1dgTVpS92D5hqLEU09bLSmfqrcwmhEh
N+RF2P2EfcYthH0VtVT3VIpEvA6wpf6StMEtpLgt7FUe7tSD2n8bqeH+uX/Vuvip5n7pmw/rScq/
/Va7hTk4L84PuQkCQ5kbQ6rp/scywzwQ9dvcCTbxrFaP0DeoRdU+nwzv2UivlShtLOQWrXjk7/tw
uidoyZQMM3sJRHQo2gcAw/bdWDNB72jrC+a2eqx1YCoGjg7V3fED5v9nmR60OIewlBP8Ps2SgtzU
06jexAKw3carvc4Ijn7IYzdfXqL1Y/ZoF9NCxOykod0HhpBodkNsfDKLRmKQJcXil3Im/3u21tiy
6FHQNomf0nxlupe0Qr0v4M+u1DLVLBe7LRF0C9jyXfuNeLR/BUsVZhDggPvco/4ic3Ex7DWIXSuh
vFJbNRQFor0JNo/2YWNUodLpSEWQ95+bFzr+yPabdZPLpC+VUb2xBsFJlBsWPknfbtsfw76tRNiF
OW40Brr9S/owcAUAKIrKMRmA/uKcE6h2ZEBe0Wq0ShAYb0Zu2DZK0XBBPk//YuwxQKG7UumphPKc
3jMa2opP3C22ESqyIgV8trVXNsp50k4TVMZt79fDWGw3ht02AasO/uD2CGKA4h90AG0tKMAn0P9h
XOdFbZZq0X0dHwraPEDsE+uyg6uOnrAADD69S7Eyd8qpaI1QUPk6ZfGn2E4eSIryoBFCpPMgCCEm
GakuouHmVkLecHiixMa8IluZkjOHCRdg+omH13+pq6rXkADT+EYs/pd7o6/g9vS7kWIIN528hTde
TcVz1KvJ4Ia79xddrpc20OTchHVsMUzKReV34CBZnPSO6tuOZ2FNKF0uOu1ozOnKPRr9IzBTlkb4
rlx8TANAHciJDgqVYDlyFNSUMoQAWtzyVf+mPvWzkET5MRx3WW/szqnTM6NgmPQweT0vpCv1Vkpu
ji+lUnG4qgyslEOrRoPh66gX+gMHhZcFkQ0sqGiBSKsi3GCqNcHR8O6rkv/CPJ4s1yqmZyznWV/P
PzjU8Cc6FzJheZ6GMlEho9qQ/RDPDEzTwZ1iCL9O3r3dTn1Go9juXKcegadXFxa2uo7Pti8Bdqwj
ZTefLfR8/jeLuDS4dcO2qxJQJq7yypndI3IZDSeZOhPvdVwn7ehTh8AaamsE2g4K7fkCYpqETEf1
VvmhanmD9i1PI7xCYz8P2IauFGEm0hZ5+u0uzWVkO1ZYk6UEYGL5iQ80VksGa3D45yZs4SVdu+Wg
D3GCLmYwe8Y7+kPT+2eLbnPgO5cTdcnRT9AvzLQI5a+lFBf3lF2uvFe0jhWvnLPuUVDxBekpTGp5
ebaR4RtmSZa19NaIY05l6/o3Ebt1WmB2zYtDDDRECVZPiAOLdvV4U4Ts89gYWZD185tcmFgdH8oH
BDT5HaNb0CACfm0IJfhs+RJwFrU4wOdptybT6yaQTKBMVg9SxGOe2laCA5Y2i0SUkCYgpwvDYfns
sJ0jdGvnZxkPqwQtBH2C6FvIKddB0m6BJyxfVUZaNq2WBHN20Mai6DWnIfzHY2vULcBFoTA4eOOp
YofCqn4KC+C1omoaqatw22arUllYGaFL1KQScOKlodptrhFNc20gY2sIFvlmglVqtHkQrxN6SVG0
arT6ohoLWBRvr4XAuNllln9f6LEUUFkfutCMuAWDbeOVV5eSEzgRPfmUkavm5fze1EoB6s0fWcVv
U7h/q2I93Q9LUeB8i/43WLngYcsb6VxOG714Hv8V1W4gNeugBRN1L0t6egna0MP5wVVA6NxKQvQJ
Cuv4zoh0q/VG+LmT48k6yz3nb9Z12ZhKiqoBhSqFRPp1yNAIBgH7c7DVYoP9h4uRe0WBQE5h1Xkq
9fKyytHKzVAEmI5rNLx48ciTipmQn/SRI7SbVlMdAVWGAMAT4jvGXYqt4figjT+9wkODVvg/MZ2+
62FiM65Cqn3ZO3oEnmg9HyqGrkDymNRzEFWgaUS++FgsTT567u07X69tbb7VUK9ioUoO35WyV7kg
m0yVaO/4KMIK4ZdmM/mEPBwJtwa1yvtUcGQ4H7SgJeG++Hf4wi5H1R6rL0ItpIcAaPOP6vUo2ooe
P4aQ/Mw6RBwUzxZy78J3yqKUb5g/OddMee+CbmxPCOwYXb55fGnnga5uOOkr2wAKd2cmJ6Btmf/W
HaIW4ufhElkFUQdoiYkc8gjOrCa3QtgM0lVJHa8a4J2yFr+xxBzjwP7z83R2z9hjp2zn+YML3YA0
U4xZ+mJZvgdIidU8Bv8HS0gLyBhcOTsu9W7W9JBTdNxyB7IcjfsHRutmtEIx3CR3hyajxycY8cxd
65V/34FWvd+2LA0pHdcqloDTHOGk1zb2fPsTxAC60GTP+dZ/dKaNGQbbiLuJoo8GaDqC7xNCtvYQ
4PlulTorWmAkeU6poE3x4v6bt2NbrlA8HdDxXkEInmjLzT/uaTq4zuLyvzwqojRspnBOr1PqQz2e
za1t2SeCBBrLzkJevwFxx9if7ft+rB13JT4agtWrFxYxwPnSV0QFwvYfZipmF8UyiJ3CmEvGSUjB
pBv9qvQvOXeQfbH/1sdc3cBHaL5oCPFVNCnnutrrkbdYYdHsRKn60fjcStD2ObOIyvQg/AD1zuQD
GpW2lXdTeuNM1AlPseAPf2QUeS3DqIwZ+eVYhIqhNwmpG9B4EkX3J/YIKSz6lqJ+lePC9LtIRcoz
Z/nhkBpfWG4yzeGMg5ZjpDRvhKMmVKhHH0SkgY8pbb91VewYU/TJB/xtenCYukcpfaz/Z00OplmR
E5VK+fOMKsQgK2QLynG0k33p0OjqXYentHduVfPT50lMb0IJhuvb+EEwxM+Vp7bMxUrbW/bv53Uo
EXJ7FDIKstYWaHeSCed2MMQVZ13Ite0+GrKsSJ2+CsklhubUyOOL2wOB5kMjntdSYFhRIjGbfAXl
jraa0ijVtr1ljG5xywA78U8A9/VhOQBbJ8MFuQAJSFr2hzvZZDRjnP475IBjgBm4KmHkbHgQDzK9
0/JLloS9EWWFcYGLzFg8zvZh+Rn26C2QynsbxTfsm+nTAl2HYRme1z18JKUMsyYD4uhk4iN2bIER
dL3d4KC70lWw4x3vqcnCYFhoPheuLI8dLDUlU5+tHW8t5yBrzxbm+5CaD+7I8DzKm8trYkF/DXIK
fMqgNDtJUuJdF/2Upq5IGaHjETNgG6V0mme3gg5MygwLc9X62SCriX4KRFQj6oWJciDWT3a2ySIS
9Iplmr+n4HBoIlY1sTSCK4+6muj1v7JnF9o6ATS33DlWpmPD0rXP/3eYFgXrRGtiMHrlWrHTKEro
nT69gW+NCo4F47seehEmAga5/JhkTj8Nph4F4XsPWyMtpx7KGltdwyFhk6ZtWAan5wgDn+lY9sRh
7FNxonI3rqY0AMh9HITU7Gd7Y+0rUro2ICasIhz7V0WE1nCOoWu4R04Z6HSPneH7pCHlFmu3RTJ2
/Cm7ogH3Uq5j5AhjqHx7n1PR6HGkFbR7kdA84fDcoYF2VXDry3PDbxWpb7WhiKI0g+w958dqhaCP
KlDXdFZVCTKZehEXeGY0pA6ddYMnbht6nwxJxgcOEAV05NE6E5l3zqcb1PVpAsscbjxiDS3ik8YS
NuggLq4O9qHxKXHlJOV+IoqNso0e3kAauKDCaNANr3h+RjXnzqitRNh985Yj8zNW3uAzTmBs6MSj
tAFXDxL1OTUkrdG4CHVFgnDo03KiEDUygFJmMAZ0S+f8B5Eg+KUjQ4L2xa42H6RaiDjzLIKEpk9V
CkC+mwT3QlHbuOCVXtb2MeQ4PTsLMStZSYRU9xKbLV70xFUyFNREPVD+hg+XUVcx8LKgFtaGrB+W
4dotaiMP9hbVGdOrwKT3sIBfsqzErqzAYiQ99VJU+4I5wE0uRQMLKEbDsCt6GInNlZsFkZTy+WbL
KMzM+MeunQhp58dLrCC63z2IxfDS/g06t8HFplJTaMbuPnmrgmBaeBXFbaSVomUvC9/mOMy4IpV+
7t41d6vGIddYgJoXT2e9sCSMy8neGElCYMO853XErB8xtOrBdk0Ou6emE8n9/0oybsRkqa45Zh+9
uYm3Z6gBWjFjoyorWAr9FzBQCiudOGDn7CnCF194K/NdugXwFyK09tuAYptW6DRbpamFCpZKpYOr
Hijw0iFhqp2Dv9TnC9xQ4xcUF3GkrjAnvYPkEs4fPS1iZXBAiUlhQ9VN6g34A9T3qi4fXICOrvwg
RsEYYH1GjifKOme+4ZkCHMyXib9c13O0aGd4QFamkr/+HQiNPzYAeGE+U3sPxqO1otpsP+She+An
glVYWgM731IdRjYcuxMFdgPTOdVaKcRxH9IzJUCflDar89BB3NOyiFb5sp/ciGR/jWx7MqIXN/IK
2s5Yu7jxgrJMWwepuiR7anlDwbg6xq6OrbS6CctLjhS+y/izVjGuCzmVZDopDJyziXwUQoljA7eG
xIGkrkTVJmCEt7mD3ri+nAYrM9ICOW0SM4/BRqkLWHxPejbYpQ1JoqagNPtWuUYu1oJOcZQHkVXO
xsGa7+T1cUr3WQtQ0YpbY1ecfyBxD58xtdquWiKzVVn+4raDfttAXgaLQTr4L0uuflp25Ta1XfeU
hK1ZZ5MLX1ZnyYbrZv8ZLmMVTsn6TKaBpmz7R6JA79ZmoiFNfzNzBZfnREsF2t7EEzG5ZsC1O8hM
//IvK03a3qEolcz3TsnFwXnY+eIuRF1ysuBp6WR4AmArjvmUx3UMCzpidK3py+9QKu6mQCVkAS03
xjkCb1gg580Z9WslrlpuNkQyJ1BzfAvxztRq4J3d7c/6TfCL6QhdLye+R+NH5cRXYdIO8MynLEnk
8fh94J40z6jLoOiAXgSn1EOvsHnJcmY0Dio7ZxsDg+W9113ipSe6vxviDKxrNfhQ5nRlKB6lKrF0
+Tlo/t/HufesR61WTAw7I3xltLj2B5/InCtIN1/1bjK/M8MWP9jx/lzoLIVl1DuN+GfDLJzFYJvi
etxsl8C3gaBO/Ng75N9Gb++hhMwr+GVNya1WIbNnj1RwI5BTvp/IQXTIcrfE7YQg+2J4a0qO3RAf
0NkXLqyfUv0Wd+oUy8Uw95KRQi1AqHpgDWSj3lKoL/aKt0RjgR7oW+wymfbVV0DLgapuXZADEp/f
qOXY1jvJyqydumP9mKNe0CtoqCGM448hW88kR8iM8yoPMFgdyAK04C3uxhqi4LeoLWuSVZX2ytaA
rwqpUYo/9cslXW4K6QFxRId8gyIh4nEDXhzr/Y9vtC7JrSxl0J2tGKMmIRJWWeKBvHcQhWm0rVGG
mGKg65ItU00UxyQWChMJkpQnfKQFPVXW8tC8gn9ez0WwxNRp6onMs6ECk/qMw44fK9BeTbN1vqSX
V9nh5sNoXmcGDdlF/ppo2Eg634Ionj2L9+ZwP+PFhanQ0m1wvekILPBj/nICarmQoMzcZpp4cmlN
cgderij4AhPAXXv3d7imhMaM4wnZ+xPERAfncSwMQfwYPL8oy6wx4RpcYV9jrM8FpWLZEgBkd7Fh
PKYUcVSPonHjDOX1jI6yQ0VPY3UetWmZWohEh2wodygGHrrzYIKJ/y3g+JlU9Zt1WZzuxBx6/X5d
2aPVBFwb+RlrSNnSUHKDMQbRDf/7COsgcc24r8ns01QJZzlMHMTzWTehuhYP3tAFvmkoFSFFKWCp
7PS3oBbVzGycV02e5TvVYSImmW87lEdzslTcQ22yPqZWQY9d2RDzhT2Wv9nu5P2fJB1eSSA2gRxe
D3CTfE7zVJ/PaF+7SsosmZCNuHnp/JVeN8lPnYnUBsdLDGw2onygaAO4JPNgmq0ulMDhv5yt5JkW
bbejFupjZAU4s8JFg78SLB6d2jDm/YWW0HObu5nYvDJQbV/aHLQeKrU/le+3u76naPYU6DKC778G
BalVPkLF+7VUVC1lfQhEXQmUe+uKG0ZLNVp93bRUB6rHMAtV0Ic/l0yswQCdASFCqSt2A/ipDd5W
xoqLg6Y/Xm4TTJ0MGpVieDWvpMOpOxEVmJhA1R95QKD+E7jcQ094c6DqlU46TnW0FwMdGJQMdNC+
IpgG1uMJG/vwbXRAU4Zag/PKRd25MgNZuUoVoUSSswt6IvmdasfE/8DAki2vLgatCmNK284WQMWt
9uySUqNSAsBigObykft1xui077p+t7AqnnOosrRsXXoIgIGXhhtMd27o4/QnZbf0t98ye99k1NlS
todFg+FqnYBop9p1sMD+uS3/ZSbaN3Qy3ZK9GVVcr8SRVhrSZjJxcQYQIvrNDHrK5p+1kglQqMYk
029JJ/Ksoe1yglcpXM9+vLTKdzphcXZdjdIx5upwfLHRiavcY0VgL7ZAcIQCB5k3aFX1HF1mI4yO
FgBMKIWwGd9fYVqriO58hl98KogtuTKIkyWCMCgPhy1GzvE/QdXtzl1gK0r+cKuAj69Y+EWfAxUI
B4mGYMkTRoouxDzLsVEFSTlViyO3fDN21qCPjg/k3AUg8e+jzHF7cXvRmueOr8WK4ZFDIQnyz+81
W6j1n3O7EHLXZ49txn2Z2WOiNeWd+2vHpLaQbRfvTfHf4q2QThei/Br/ZmaIK9B8TSQ6Kx6j6xkK
2GpR/OZ8DaLLM448SkpokRO7vg8os3rR3OjQE9FIGnzdNynwbPBWtrNtqkm8/7TrJ/9VuC+fNlp7
0hzLK6/cabGhiYoHjmJDYJJSeFLUYkQUnIyAHcaC98LFIm2NAvmQGChGYvSfUbU2kywiWFC8pCV4
9ohm1yYvs8G/tS3nWiprfwXQRwsSb7yuQjjhiOWQVwJ7XA66nb9ahYiQys50pJ5hiXK4dEEsw8UL
7UlUE+bfdY88aqe+fNiqHiDfM/s8kUp7caOq4gcCRItMleIvZy2DOumgudC6nRHoy7Fjl+GMalr9
VPVVxdmzOwPw5BZnlHnaO7fR29ShvTMWzuwuNYDqFgV/bkzdFcJn355dtRmOpNK4UHtB9lFX5j15
uuc/X1ksHCHS5KR7hIZ5XaB4FkI5fwIksfh1b/hepqQQYhXWlDWL7jr9OopW4lfI9sewIvZd/liP
JOXnbNsHMhvPImInuKbfloFpYvzQmLfBqQxz5meDsBeOUplZBpvlRI+93edpqZM8eff12kcPDy6f
SDkG1Y/YGRUeTL6zR3baE4xLomp8XIfEHMSoA3WGdUl3BpRkycFe3WsLGSKAJpyaSbxARe0LrJR/
ROqNHvGH/luTiVXYC0PehrPjaP9lvN9bWh+hiCOsvsvNEGprbQ4K3wIpoEpdur3f6sZTiMKzjQXD
aZhdpxlwpAEkkWU8AJVlYe5/ZuN6J+gbZTq+9jAZcj59qjerqfWIvSbHocSmmLQyFd4JkfQGRX7a
vvCD1OP83ToqrO/e3ujaOQKN6yJNexx8q5vHY2LpRRqhQjj6Ap57icmfGPu90CeHy+CJ4/bITeI5
yr3SXLtfcFdwxk/Gj0fOg7aY5aFTBU66pm6vXLzrQAdO0/jQHNuO0zO0BGKt/MHGQejvw1ac+vwn
8Iaks2j7xwrdpb7oCjUTLXYxrvLCeqU8dfrCCS3LZ/k4WRfsb8GExBfETt5kXmZUWNByTO2mEmXY
nZpy3v5GRFN0tQIKAHt2RttWtgqGcytybzeWAXbrUDlAJZgG+RGMRKHR4Nh1cB19EIddAYWfD7N8
I9nnw1KzfWjLX8gFO2omSnIYQhAvBsxnaEUu6Ig9lc5iEE05x2YPIrfjFNw31TtH+uIyPglD874k
VaDe16d4qEUyZ1LpvWom/vKwfqdleFNptbMnduHahzQgE1BVuFvqQ3SS4iP6qbBbjuGI1SgDn5KV
Wy3da1OAE9Gi1VYgP/d56Uq+TlsAso/qrZ1i8/Z2wTyN/7RDClRXBTVk1gZ3K9XDwhCi45gPsxzB
HPJ8y+UnE9e5pcmAr/5c9CbF+sZmktxiwF5GkIKJ6EnnUphsFAJgCdfzd704C02/2hINZ7ulK6WJ
dtp9FbT9nPtKETXgxQWmVfF48s6BolGmBs9TeuIGICOhrcpOwf6wubTFjZFf5VYvQcLPQ3fKKGk9
nd/eYuELue1j0E/OcCbq8q1tvnUr6M8T35s/j6h02PQYIsYj/HB2pkHKkVVEe6oy2ELGdkl9QdVZ
nALrrZ79+/TD8/2GbYjHpbqFP1Lpi6yCMrRiEg4PEMWt/p/30mikc4WSjWHllZDfn0b5CusqepPJ
Qa/iSEqFh34I2y2i0Yge8q68HkUlSkZrEfjT2vG7xAEJeTQo6ebsBpMaOlRp+wzYyOfeLfVYK0E8
r1CqyUDSCHgX3ZHfA1QoFlELQMeB8o/iP0BKoNHEgo1Ml1gSjr8lw6B+7jrG5MNz911jRK/yZ2Ik
FNUniKk6YYYr7IY6rmP1/KLIxCAjn6txUjTd6D66dWkT8axZ56fos0xlicIxnMdKe0o/FFDmAKu5
RITwzvaPDifPxQU/wmT9HE/LXtoQ5GaXV4ltDeQXY3iVjpWX+IH7g7XjDMr3Bfc6YIaqK4WIJzNG
B1lwje6xKP9tmYlNX8yn7MnO/efwazcjdSf4n2vo4LrOyggR5W6Zvir+iVxiUbguL/FovmcyEaxU
r27M4djETB5QKww5wvTi6EjYaMiDLA4dnQHKWIFixGK+ZkyZmMWX1QchyjqP7qLC0dqGHDe4rVu5
UDZnEzP5V7T+nVCnMglJmJdE1QqbGjvGUqhPzHPtXEAbcOmu9QaLDCiZVqzxYnUKrheiiSQxRvdG
JVpME2BxHDRbimwt+219b3divBfHT3pN5v1bQ4GUDP+qZ/1zD+DTbvAyvAzj/roIbGXDkqmvbMHB
ZLZBQb2/josVvh7zFHX6VD6vnfwlGVyp6R73p+qH5a9cG8nh3iLqMIpnjOs/JgiKRxvJ+em9Tc5h
hpPCTYRbd2+IeZRK1S9p8CMHOXrZchq7ZbvnEcxvEyREAVEqsuzGXPZvO2rydauJbEmId7kZnSZP
+N0WvsH0bKFYY1zpPgLunzNlemnlnmI/99o8XowyIZTI1hDNuCOK7ckbLiVH8/lO3ReViIijI7YM
xKowjilZsCQEH9zvOwy4OesrkZJaQZuxBvZP1caZHVln0K+dlPIP/ogRN8dGaOkOQXPhGL+ywkw+
XB1c+NwUkFdMMfOi1aJkj8EgCd7fCFWL8DVi/feavFsHf4tyyvpHTH8Dp1995dq5sbmER7lERsaB
Ts43lvRMGANkKc0Sz6pkaxrNQM2hTA19GGAHWfabrLNqiKcxM3M7QLiqy3KPIVeNAEbMIhBNVURW
3QLpfyY0XJ79z8+oMwQHahYj7Se6A650MRN5eG83soIh9XSYgR/4TwdzgaFKLw7n8goteVcPRuUA
QYFMhFucSyzWo2fka3VlUJB/D++wlCyHIAJCKT9mI1IR1GfdP1ATPYcyE+QFIbwFIwubCZGFCJtX
vjxEGcK41MtxL4MbwQyAk+IiG4e7aHbl641szlPmB0ZWi5ZDuLxNSKhe/EozRaG2H43IoC3Q6kRw
DYm7vlvQ1Vnfkf5RbDdtGMND001yYY407jcPBwNLQ6lSTW0cJO1HiCNiWUnf8RAkLi5vK1BnMtYz
5Xx/ByBIUfWyUNNKE2HSOxr5uVltXp0tYB0WvFQWCwcPvg2yPFIwN9dRUi85UwFSJQjJmesH+pOI
citbHe9I74ROoy6RhS9OzD0N3ro/Lxfl2KNd/jf12kUBAddh2Eb+RvmKN4zKXOTiJLVgOdr7hhJQ
osuCoozkJCQaVcLNAO3V3ejZcuNzUz4tzsmH7a47h4HDTS0lZbVrMUhjVIb4+26bIwSVu0+yW3H9
9xXA5VPUM4pBpYvd6ZKquLr41xURP9m9pdOsZFcImN38wBq9SgoE/PgQJ/ALXkvq4LXNKcUpbhHq
QE9nAxbAa9cG203usMvlyKNK3595+sID30vpPzhHqk1D4XgUHbuOT4ax88Ntwo819dVs6gDFMPrC
TqCD2w1VI6TLJ9ywlkhzh+RkToUsty4x693SkigYJnsqMxXLKvtHxVQEn82b43qbTwgzXKSx2lV6
PvKvpII/bzsCrgW2P4QTra/Kn2JRCR9X1EG6zZe2egSf0NdNgLuZoeHkbXIKH4F32iRCuqCIh42l
rZwKRYgpUdSVAD3zAesTwcPNRAhCudwCKcFZ6MxRyeRVMklxT0ZtUPbhTx2eEwJtEvljHy++rK+s
ShgYeOJmonyX8wiyNQVpjBcZTOKLDjEmjHlN3NR2ecbJfDF9SEnP86j7DBHpoOtnl03EHdOQfOds
9juYE7QCrMWSQLpVh2TXT1UDw7GxgqEXF8OeRMal6VoNmb34TCH37HVhxWs+c3myTqcfsELieYfv
+fq5n7VV3qOhK+FK0N04rzWhC8+pdb1/HeorFLW0TEnlNcus7SIgjNUl/2fMV/rgGZn+PdWa20aA
GVz1RL/Mgfp5Qs8dWauSe5pm9QQ0LK6Xps/t2DmPbQB5kI1vRNJe3L8ceScn36hVPR6I0tKrCggU
jhBaTvpYWSjQ+cVF9rDWxOdDMwEG32iY+WdlkJBLLKVA4cJ7e5BCjLdN1ysvDaki8Carfn+sVULO
PCnhgShlGa1UUvXIDJrhIu6M7gSHxEX375TeC9hvPEH5SKOlLUprFo2TvPp30KUYmE3dJviHWrHZ
2bA6TXuqMqd8DCG9Z/knGwoTI9lkTQFowEseUxdL7FBK4OcW+U+cqSqoEm9ehnFJ4aMKUVjqy102
YBpH75ZxqxFkL8sN5cmDTUrOWUwrtusfVIP4nGrbknXRRzbvixUEaZkQVMfInwVwz1cE9osvvD5y
v0L7Tjj/SaaV9Rg+Ib6+gnoJX5ciZngNMKjWrIKaPnxvgSFY4jravQwgy/fuBLV7S5LqiZhQbePv
RkygGmsKGJ+h7ioP18ZRpfldBbUFPuYUD4NQG/+G6f6e/tlKojIQRyP4oIpKEUt1xzHuhR4OkFQh
Mte+ST31lrdtjOFrGjnrJuGQ4a08ldFLVA3zrMpdIRMde5Zm6hcAdvbUDmFzV74uy0MhTjCAoDxP
Arm4y/qnVfCZYgcemxvyvAfTHhbLJaQac06bVzCMyQlTheI3RMT0o+kYUp7ryKxDmY0KAe1IfbG7
z2GJV0hw/Sd9ohl1tJf8bVhCaskbe8ln4PXpPYuMoHjaCjI8ZSY9Q9nj0IekH32iWs/fHUTAM5ra
aPq4DXhk9aKHiqoOkVjOqt7eJJaq6swFRZGCLnuXpPj2YhesQJ4psFBLglReg0QJWrRTDJ1tv2mS
PFAuIBaGJHl/vwGh25xfTe9LAqDTCnaKo3mXWxbnr8mcx0MSAd3ARKFtSVMnphbyhKmmiiTgDfGJ
PSBvrt6LSgeao+SOvcO6y9qZczd5+cnW+bIo8QWxPXH4EBObJfDoepiYNmJu6BSEZoISz9bOvXif
RqQlmglsnaJPB2Bz0fvRDMFEaBvPUIWQMgc8J/jVppxX8ETk/oZjFzD4/LaH6MAN2eC4Kg8EK4Xx
Q/42wE+3CRdm5JlCLbLYIMTo7Q/0dADELqbIFixA2c80kIa5f9ApyySeWTDhAz236mkGcap5i0Mv
ttXf0ohJ57CRKYJolHJdbYKN48ivYipD3WnewQj6xYwZajtpuVg4Vp55OQbLZkbYkFYlR4eCry56
o1G0iXtyZAxXu8nBk+9dlkIhLH/P7otDBlCUt9x3qZ2wgWvoJOFWkCJ8JPuAHRMsnDY5GZHZO6XS
FwUIR2BJkB9GhDcJm/r598+wExqz83or+OqHIH4SpG/Dpo0zqH/c88dKxrO0hMExfTPrnAeH2C4J
IE2mHOPxg92WWR3Sal1uM1XaJQcZh7OXy60Jo7oyt0ro6Bae60PDjlkCjzP6DOBy8nKeYbCSkhme
g79qhFX9b2205jIfDkKK0Q+EuIHNpEY1JSBBCBsHZ1La/2rYRmlG5RX0XAnGnZ4knScT6FeCWUnI
xamVjzz9sETYMZSMvFD1e1fAXENpYfpiFIwF3ZSqO99Ci4IxLyaOJ7Va8O9kUS3GCi65ZpnOa73+
1COIrTSpDzA9/4/U/CvdOhSONHoZerYacWcHm9BxM5oRuCHmLQYa7fwSO1VJnpeCCqZh7nLT4V0u
gS7VVsb2C8X5fNwGJlPYxRjBggiBFK6khwssymLcbAVDk0PIiz5/zPlU6LrIwCFR1f8NYnxnTMpK
a1TyTnTAaw46xwnObQiHbKCWD7giFhy784HFi0mNE0ydX0kic4F/3Q+tOB7x+sX9CDfCzUAekKlo
9cFvcgqu2CqeOqJFl+TMxqYRVIYNfzsHwJfyiJnG5eej7kjrf11vJ7Kk4opPIeM1aQ2UOImqBC4d
RvYaC6gbK04ra/tGH7diosM7GYMFYt18vqsWq4dMQXnSkpH2whB4QOCBVbRtxTvBVCS/EQHKz9UZ
kxOGs4dkhsNIKkwQMfHevyMN6uku5qAQ4g/DsouNSiKxqT34JYFDSnGlCd2z0TpQd5Jthadb7Ikp
VIkNfnn9o7l6QyW+bSzndDilc+45EJiGq8JfO/bGB3hbxAaWWjqmOTCsahrwsPnIt69Neut5wpWW
uUp7LNlZFLStt8CG6t5UvdW27OHHyazwrNQBCzDaE3udlaWicui3OjyTXD3CHY8lIs66xsxW9G5z
5vsA06PP4ZjYKQE/0IV8hbrVSCubK0ypV2fgY95a/zT0fX0Of2pZjeLLgFggTc59AWzkLjjUuEQS
/dk/pATOiAaFPcvWUv1nxJv11KdSvNi/6poJ9KeGA6pYxWJ+4ReD/JSGhydt9RdsRLg7QVcypIGA
hXjdYGxZEpfglBWQ1ZgpApmOZhBFeh2ScYXD08VCbj4kAL4jMS6E6UN6Mk586u/HFlH3ba8Ktg6+
+nfMWDYSR0GKEe/hhHzqYKPcH+ePdhpGKdCgbcy7EF2V7uGhCca9TttWFNOtsBvWAAviJGick8a/
0PYKGwyITPthfqNkQ+IVNWZjp1MnqhrXL6R+1s2IW0/tKbe4DdJKoC0+FlVrp3BwTnA+FpPv2lpB
nU9B44qVq4naRXijm8UGPnj5lc9BcbVRigp2IOTwdoG2jHi6OBiuMHhFWnXaPc46NECNGrY36jdW
8FvjCDw9qsH0Gdfm/gHmhzgSLoGhNc0hdwnIvD1jBH63dcLNvEHUL05/KBLbZ2g9R+fzzYATDqv8
46B60ZcijpTkDNnOsiNmr6ig2UA5/L3Ky7Eek7kfy5EDfMa7odAkCtY3fLzaQn9SdTpmfe7iaI/R
Xag2EkjKhRbTT3O1st5G/Fsun/HVffp+j/D9RZLRc7s44sGBICPDJh5gyX+SWQ5lkRRPzSctE6hy
bfbcDXtFfk0iTabZgnHJoJ7pADCGpq8Q3ZKjekoMMxtVOq8exX1CJXiVwtO44bWY98vPMLRnon4O
Eug9pBDOOnbX6y1KVec85AF7lw29UX0x+S1QCm+M3GoV4MwEifP6tKo/qxaq5Ygq+oIdrn/j1kV2
yibJAMiKXBVhOnlwoTT8WUrrPP/YSEUkoXMvpc1ON5uPgmMGldOoAlSqG0/06YatYlBd2c1Mzgiu
ovdhKD07rG3G9/ztVshVQq4P5ROAf8IzZNgtT5UpCwnIkWPLgjkZS2TKlLw968Uag8BrB7g6a/G7
DhBKRHYftGWX8soQqsHRN087lW0V8zx0wKp2DsUUwuuflIH90tTLi42dB8eAU7+yiyFZXdHdaRZa
XFCDMbGFl1WUOjOxq9vAzJQ5Vg/f9HYUL4JVqNXZRH3B+/GG6sQMv1BNQZXyxLzl3e+AJnvKrsjF
RGtOdtERbZoe/Kd0eB6Xr2RYRe0PEaCILJWo5D65BGnR+9vZ39JZTnzgnvjA2UQiggN2llhIGiUw
Dr+cOnzzaOZxkiLwdlsTu72strnRF+3ar4aKFasMsRjGPQgNticyyD4FvNCJXaN+xzQbY5brgofp
W8nfMqVUqRNPWgploPUzvvTknpaAZNvAijUTwyIiN49rD1YuK+2GNAdC6PzXXsRtcGzk5peQJk36
8wb1+dFS47a8lB8FByp4DjZughefOl5jgjKcLsLv7l+s8kGm+D8fGqUQOKJizcmqCT+w5O8xsjmz
VlLJ8rE+BK+0Vsf1/M1x2W8cgTTRmlssOO89Z5FLQ8qk8trfra3QZYIp6YIt70MqeK+mWvlYDGtq
vOub0AHFAwwDvitYBIyg5kX6z+wQXwncU8Uu0NQ7WGjoC2wdDTTHjmG6F/uy5NA53UPvePl+iDvU
M1a8dwLhplVzcowSGOe4YNhJV+pVeaX30X9w4RJvmETakD3e66razEtvyh+4iMWK+Ux44a13D+U4
fHBRbu5q6VUK18Yq9SsilTLMWJTzyYdOVW5jk7UXrwRQLImBmD3PxuiadXfjfIE+GABQDzGrxKyS
jSj9pV5PFnN+LGqbHkPIYUQEGJTt0ntDV2xWl6pAMWYK6J4+AlGMUGkV5APiCINOzzJThRo+aNUj
UYckdOMC9bJGCerMSof5C4egUFj+H9PsROwWDkaM7B9a6O86azu5hx5crZIkjDvsWnWS8/Zrdk+m
v1vzv0ocP4HHF8qbcP7zdp2UOkgS1Ah/IANO/IRN/oHvZIfXFyu4TTrxHt9tOT2fIAk214tOk+l3
5AYVzMWpP59gtb914NP+0eVSCax145E3xB8uHgWLsHr66k8UuzZ80h/R1ihri/CCwZvHMSKrtrFj
cxjJW3N4SAhnIgYknV8GsYPd8x1tSoZwM11snSQZMeekuYo56VXVA46j3EvV+v47fBTxSyTh98Ca
GJvXPEK2fzqGcegTn3c8dtn5DblE0ui4r5XPRVNak46ASBHKAtTCw6ZCOvpy1QMDv+Ln7mRJuc8P
s9Fjxn2bj41RmScQbm/lC8qECns26Q+EvFEU1MKke4x7VnBsJrPN5wxveBz9p+QRwdxvSgeJ2o/T
pDUAPL6pI0MpcKa8ztg28TBDZsGq8iAVqcXuwl7lXqCHbsbT9GenkOkCm+hFPb8UaxrKv1YOZQWq
9Mt5Qd/9exZ2Y/Q4q402UsHH2uxHoTBRRGiSdMUWaH39zCAPeiTq4y5Iw3ik3E9NzdzUCQ+mOAj7
GQAEccqSnz7ZuxRtrD9poQuDmwM/fDkwTT/NNM1bOICY6TFR7omszIXs3vlSeQdRwsadp8QGDt2Z
OnQHPfofJQ1kNYgDxIhx9mYQoegWwruPudWLoFlw48iDgCFdjIno+mwPootYwuMrl9TM9KJ2N1Se
YsTJKsXKDFfqYhejPaR5MEWR0DlCZrYXMeuqFoNLCQlRnjqF79rOUzfLlvKwpL0KEeLC2V1OT277
zaxhseIwkpT0XfjfLhyNxVnapExslyTUb1IVShuw7RhinEOgf/RUvE7TmU63nCic2s6JpYl+VVLl
UtTerN7oo2CvFVneMF5OVbGgpUQrwb5c5jXrW/axTBDNfCXTjiA02LMS2O0EDGbGVoDG9QbAX0Jq
froeOafmrEwuA0ieNsaqIqaFrvdExpgpHlkCt2piWOVUxGL1Ap8X4MlmIBJZbAoZhN2kfp1/HWPi
dWbIxMxNTvjc8BArstWR+1Wy37JLexiAyuy8OIP1TV8YB5UYrfmOs5QckO6EfYKl98hoSPpcBQch
jWRR/gdlJ5d+Qy/6E+Ced3aVPpOCZyzjb1EOU78OzHIHICyAkjGHdyH/qW2TSYdVRzYMvjZonh/l
atdWOBOVvgLE3bjryTMm2Z37y3BXRPiR2BlcxqHSM9BqDEWkHRAmXtFIPXGFLInQ8ZeBS6crPrA8
7EtUfnROP3cNRHchO5KkeZQTbMhsYeL7uRMD6FWS3Oe7qF4LYIZa1rqzUh0LA4PinA4DapGkGAdO
jLocPDS7twtRdGRuB809j324zNbH/qs2UuCfNtG2MY7fRv/GTm6DY7L0lhpTUxInSJiEeJajN2Rs
CYh3UEokeoRl+R7KoJDAKPPGlovIqjXQdtRLIEINCYpxvSP/+/uDZxQTeSw9KCMZhSqU9/jHT7ix
PreuFF3lCeOUMyxAAmOBfJOcrO5a8BPcTLRScAowqsw9MvREelkzoVMXsgz6nv511D/wkiSDx48R
o3viL25z8jumTvYhBiBjCMrKzzwcfdspykOmR46gsymehvqpAhhqZLXY9YgncC0MdYeo2B36iEi+
mgjIPbdxgts+YLHK0+it9oaZrV1PPhg3QSfcEo9YRMWMPKVgDYr4yUC0o1hjMLesqmfWI0R7JJ8V
RQkJCgTRzvDfa/alG++Ao627LZdUy4W2ryOCW34ARfmsbDGvLTFM39fyWeUbt2WEjOicnw80mVT3
huEPBlTAcoibGxvlXgEU4TJrveusn6XWAvIXESjfSqYKh8Syw7/7AFGupQMbblDYejnoAskMU9Ci
AnbP5Y9EkXOMisg0H6eitvn+ipQqbOthwtY9vbLdMbmrfoBI30vVnEr4qwXLXCK/8A+IeE7nzs+L
KdhN2jq9Aha4Z/NQ8QZmidB8yQQe2D3eSPEU0SjqE3Woxf1EfUcLJrkryIPBEdEiQtZk7FRGaPmx
jDoWm3XHTvTSo8cvkPJJWQjXomnsCM53AvqTDMQnXvf5YmwImaClC9lX/AI6CfKcEL+okxk4/OhY
/6ZH4pp4Hxb4rA43cdfpqqzgS1A0Lc88cuL8DGlbLLwcph1H5d24Q5s6AJPgr6w1ugHFKmUtJ9Hh
3afqFce67jjOiH1xBJZotOjUjIwLMpap2F9n3NEKoo9EPtUETOhNg/0bl3aLc7/XhFR1LZr5j+EX
vN7uHz+BkgDikSawqtlQrPZGMWjngSxBhVdvvJ3znbPcMkgeMugc78Pb7BMPi0VJtwZPFzJ3BRk8
yFwZjTknlBlgc25YNrvTAJj9vfeVSdFP76wG7K6bx6yhms+5fSDbc/G4/ugqE8a4UZkLIul0eorP
3/2Y1RgsH6nEMLX8YInSLaac1qNgUqP4dbNlstPIXKkv7zEqvFvY/xG8dNv3rWFG/uFlBpAwdLSi
1YljU5bRBGINgslEq+bAe4d2/0hnLwqWVB+z93MGeFEMidK0xnLCAWOka5ybaL9Z5XkHfUCwDE33
sWW/dBm2nxCiSFO4t6NTgnTYPFC9Wl4OTt7PmolXRZoZLyrMW6Zdea1aIKu1Xmza74FDk93MCzk5
DlcY29KkwGYjDz2Kua0Ds85pEtryykbkPco1JF6Ma5+Msy0hzzlVqQ5cVqfc5eZCnICFXFAKm1DK
5cc9Aljye2dj0ahRUUS/a6q+uxf56fTwTwrgcDfbCCkTyxnsFofuFi7k90bEBuWEgOL5XHrVe0Ee
nDlOHWWNMbBA0zgDnQQRQLtPPaWVD9ViVdyOwsGHG5N8tltXpGxuIP9lqXlX6bKb9ExHsFrFGM1h
0cD+SfjbievN/LD3vK1FKm2fhLE/JT7i8immLbS2Wy97TITNQmD5ZY68iHe3JVAcI/FxXzyDiqra
BX5PIMs53peNtYuOUpIocObpD3qiz+Exexf4U492OfuIRuIcGUvGmOhmQYfE22JwQ7h6bnro+MXR
WOK4lKa23jeVEGYo5PjxsBRK5jGqWp7cr2V1bxlCuwSzflE1d6rwK4MjIGN6zFbEEn4B+UZ7ES/0
HphRRLs2dcnLreL4BRo3oSxoTD3plOTbhS+fFRoYsa0TzEzp7lSnh2tB0sjm8doWsnZH0zVikilo
pJBdTwvoGRvcaGoRkGwOs+lX52CmDICAC+Xk8hgxthmTfl3clolByZW8SD6/hrWxCLwSDNpwLuwO
d0g3zLrCsvErZW2JCrk3KAXYFOdeRKM4aeUrPEE//ifb/tIEVfC7px55Ymy3AC8QZuqu3tJgJB8E
3AJ4sdeb//8rI+l3ujkHo73AzTR7q6xGvpoqVhRApnZhJEWjb9jy1O0ZBTFTIF/hnhlO7JJ00ndq
cIqza4bX4aCytBHGyw5rItz2IR9PUhfcmVP4gFYQSQ01p/2bxQ0ehUg2ObGY8C3HxFVYFBzQXzyv
R3UVelkoRvQLZx6ppNcOjvPhbd/Ba6K9ZTRkT7kL20MbSGQHsG17JY+95Dj6zJgJ07/95iksvFxK
+49+HUTJiZeLJaeVqJu3m6ZiwFoQFiOyRHuRI1ISK6hxV0Jk0luiopdPdY4IC6cMC/IY3EmJ9qh6
LYJq87XV1SrpzDL7uiRGOnP+Zd91YbTs81QcLKRUgzxrhHFod217W9Vl4VBAqoYnhLZG58FOuvJu
q77edzksW4vD5oSjlS8e4vkOF8Ankow/om5YwiethsdLsBv5oO6JONGiLBPdezqKD9CA66bONFyH
AHgyVSftKu356Wvz3Rym0C2P2ISRFheGYIbf3VxWIqZd2Ipo/FHFAAItQT0CEQk74K154AkkbQsM
fLvcX0JDXJh9J8gYuaZG1BcmcrAO8iZs68CAIknb8db6w3HzyhleVvI5z4SJcmaWGQGnPYZhTkG5
qNrmiv68fuUEx6bp6rLO0ErFEkfPvLmjTDQ9AeDTMNmjpdpzLuDPniAzZCE/Ds55T3cYPup6vRZM
UxVquhodJzlXEX+ipjwkL6zBtSWv5dqc4mnXOLr1gWWu3LcLNnxxeJjnrkvRZQup6QLYzNCYf7e2
iWMXwpRyhvp4C7Sb9FiDu762Sak4JxuRO/PbgzRFrkvdsKeGy9t0XkgA858WsnefGUL9+N6xeLt/
bcQW1Ou/C8KT7+06+vYBrDPAzI5giICO+xYOICsyooivxsen5lIGu14IxR/NqYkbtUJasfMwsqDz
7HJ7qqyxGng4SeB/XZ3X0PmARkxDSbcztO+ONwdpu6kiithDuAkl7Rix3hDFiPCPFDfX/udQ+Uir
MNJYOX3I6NJ0w7I+wZ7S7MKQO1tO2W0qwN8RMgrBIzBANStj3/njL574Uz0Rp9f6y0cVoiZSu5Kn
fA6AoKWIf21wqmLvfXPNhDs7PS8rVWCwElgJ9vNmxhRFHqPrMsrMSG4TXXKTVp1J5aeu5Ceju3Gj
q9Xgbmlg+e2Uj8XQlbpwaUznPpGMZcdfQsnUuOTwZDqP12dofPz1iQ1J7MweEkZ19zmFUMbchHZs
J3HaMPjxvwH3XLiMIDZrbKUq0JKXbaRE62uJATFBBwdbgjQnM1+o0aJm8XCk2/3ralFd94w+9e0A
u1VEbFna6htuc+axMrZfazf3T6WyEvfFaTA6uKx9wn0+Dk/xQTv/O8xSz39Z/IEoS+tiqaMZgQUz
unutSV46/SrgTqW29XrtgDC6IPIEctoqp7RpM6J+3TKHAdHUl2KO99/jvHFh8yFd/DsuKYLBvSVo
XwdoIccRKgmRtibVSpBqeoNRmljwysMvvu9E5LVOz34cxH3nO+j8bu+03VXpUOWtPTo5SZYt/hOZ
TRIU2Hsl3iDQD0UgYH1rnZtAGYuy8CvfoO4SN+H4SSA0dnfge0NVohDreKhS8zyjjrNozEKnvCP8
HBReORn6BC/LYoAPWlyLH40GZ8KCrcZAWKc6QU2YtbfPg2mB3sIjzzCVeGnIft0Ud1jmLM6b5UN2
ZNBKRET/HNiRQgZsO57CXhMBYrwjbiT9CaGTLQUyW2dXYQfDNO0n27IrIOLfDFVtLbCiFMvJucxP
mPkh3KFAd5Pj4HempHvSp2fpMMJiiuRuc1RDR/L5ekH+jEsZxgWNFWTc0J9OMrzZEuYBVClY8X3W
cp6JVEY3zDd5+udl3QX2QYAfq+PNyi1rg7y8owRn1EA3FYjA47BwvM7zhfR+x6DfKYMao7mzXtyl
uUSD7/XITvaf7fPU05/LYBmYZ4Uf6EN97hmB6Ame7XkDiMCYnvDCnBnrjhqa5VIsTH9Ohrq6R5Jh
m2NvN2E+nuoMB9Nw9hJJ+gQmLNxhqeh9fTLasC7RIJOoqqIz2A+vWpy2GPjTxKla/bwAzdthXIvG
JAmP2S0yVDcK42T9jUaxov2muSJCDKZJH+Dy6JT2HSilv26xRDiU06rFO5vSxoOyk1P5RjqV24lK
5z6/hbA/p68tdOQsp2XW5UQYahLjaAANjMsp0sA/UopsRcc8mkNGtmFedC2WiR/CD1xDbrsAA8E6
gNON/s9wpPDoJxp2f/822eWByipnsNJgZ0GHqAolhxtyJy7YDvqTILj+q6KZDWLPHbz6s7BA5nAh
ruZtUYkANUApuCldnLinQj9pLNWwGDTBbwBuL52I0wWyLLKteFwvlCAs/b/AJKb7LxrZhucimu7f
Ow97WOW/Kw0i3QbTGAd2lI5rljeB8GeNOEVV5dlX7o5kwvst5WR5ETgqij3VyokzLoOTDgKXxp2B
nq76RFJZ/5wB4HqWfRWj0UKgCNekRg3dXwGtnF5MSvwDLZp2z8iREsdCNIsIMjZaVlub4KYaqucy
5cxMvV4rFssZ3rVlJyJ6BD4DwwpqCKuVzaTL+Eb/XcM06Hxyw7fUW4mpmkWiCMlt7wflExogXrSV
gVkumCXxmPZTxnJ2wjquUhNW8cz9Uxgm8S9TYwDrHTybfE+vGuQ1RAqavdkJb04Ap/HlqyE89p6u
gUpYC5ksLJMi/V5322uZZ4Mj75aXlER3LZDOex3ZCBEMZHi11zofuB19C6SfOE/hBJdjW1aBSPjC
NZm696bKfbkiJvMTZJngXfvGz3zdkolX7vesyzrP1VioBw66VZ7giD6UU4P9JqY21NM/ahnECAFN
peUcKJEjWeD8aIfIu4O5vHEv8DXp3OOPww7lra9AwiVpWFIFBRy870kBfWomQovcv2I9xTbpa7xI
CaKeYsutyFrqbi5KK0KA79qAhsutLrU+ZZvQeAWV5/7hmk0UBDsZGa8aJfTCsK+4fMzUuSrdHa6G
zUqNq+lN6GMj24lB8be3wAcG8gEGsUZHxdmV29fHPpWXUyV7MQJlrjDXmlU0AZVjDQVRkw0rkCbJ
IEhtTWnDxY+57QjRc718WzBTFlfT3JbXnCUSt8SjD7Fh9HBkIxdjuOSvfwW2lFYcxKChMiD+Wpj9
8QjNHFyuLRhN/OCbxE/xDKXGfZedPVjqC+oKQUi1sbbZJaaUNQr1HIQSt22bzWIWTcCivw+Zljsp
o1yunF17TWLV2RMsS0cXl1WWALIWmPbFkC//ItmZystfC77ryvwbRXrqigQVZL6iLRXCAPcKmlDP
Z35LMqsavD+uy8akZp80WwCjVaE503MTlUoQ2PYhuo4u5JTnnF1sie6MR3vjGQ6sTo5dH1Za7VOI
C8nB3zkpU/pndUAAu8iilNwTI/E4mZ7Wz+RV4Hh6fzMifdJ+3Q1XUJEsD+JuzafkkpG5pKEpMxAm
P1eRlmEihT6bg4QOx9I8gLzay7ipEsfV9d0XPxy7O04vsDihyWyG1TiNmlZmbayGYVEdCWkZb4Sx
3DM9GusCZrOWXiT3TGjg29K+caj/JaH4zulyu4WUjE0rF7o9V1n5ooaM2TuNvBtNuOTHVUP61Be7
qyHRqrUbkhE/FhHVuty3yd3vy/28HMwXbUmmeV1D7a7ItaZTfFoHZMWIc7iFWlE3CdUi/x1OYR6V
um8rRoZwrjszDKjVNBBYqyYWmDYQZ+tyz/AOhYnutq5nc9skM00n85sVHr1iH43MACplrgqvr5im
zmDx0ypkVneeRd3z1SoE7sMVBqluL9taMvPBbhwsbDUcnLsUQqGilvwkssdXGAiZoWNqHpuA50EG
62hXaFsc+RLkmPIQqakFcewLVTIsUgv1pZ5p/sxhRwQ8ehgtApGDAqrbega/HK/2VicCLmlMiNhF
z/lCfy2a8MsBo33eAgt+kvW0L+LLG84cJTVhdWZBwkuz08siuz5cJIU6YyUqIK4+jg6fv5NXPXxj
r0vCJ9mb0f8kdQnws1q+kGcqoU+Urz/Kgfzx0iKFnx9Qa8KQ1wQw+vdimDuxop2ICIOYucCrc7Nt
ofrWZKA5e3QWATHR363KA052Togdrx8IOwB3X1WT7Ml9iGV9/1s3ntPN69n7HpnFtrgToU7F/o2M
75mCWURcU2ZXo5eeVnpqVMa+PzW1FNiNzS7goqcNaohdh3NR2KBf0QMpIrGJJBI0u6CDef8ENIc4
VtgrdSs8QuLuJBzUHlYWeKYOr+1j769AtFLajK2E7BtBmaI2AJ0AjP3q/u1lYoG/7D+De3nGyQ20
lfG0BSOz6Bu+XMjfJdVyV2xnBKohMoz5hFHxMCaYJENPhODVaxjXpfKu56Glj9XeT/V9naffRkbf
Yvzi2Yeq8t6tpVQOVJC9Z6Cpyu5ki1WntNVLRHX/qWjl6IX5CdJuPNOIa6agX26fOxK9gdPmegJ1
rZyfmfLvtv9BcFOEFqWFKfPQ9ZoA7fo7zsKqS0IxxIYC0+X0pK9uckqOFZrHnG+5vx/+oN6s/hyF
lePAOAkamHrkYNvJbbusWIz3rYEdmaDuyNGNtvsJfVLony4ft3MP3BoMMr3DNDczQH2kds2X1Xzl
Odnz/A1SOHiih+b5KBAXnnUCakuaGddNxH0TVq70krT1B/CMHU3VJe8o8ruJOXbC4Xgji3zpfXHt
JEZRVTnM5kHvX7/0ZJi+tIarNTRhGqZOqf7E7DBuKepTs9YaRCYGvFtYacoJgqKReOFIogR1kyQ+
I2d3jAqKilItO8VPaJwz9bY9aZTLLKieu8asBp70w6D242mZASlZ5dATk25dbfrSeW5naJk0JG1W
x+smZNfSfeO9+XorwrFxABUiHh4jA/O74ZoeIifYNRytCYxrMAVUoKgTqJfGiILuG2Y0Xt1hASS3
6yVt6lt/pb+69iP3sUWGkFaEfPHlafV93C4U/aHWCB5DBDzJOu+B+0XUgDgyuIawLyoYjMJSAIh3
WnfaZl98MfURhit3lfb6qp1CCzwpu4mw5KTIrZs1ET+ZihWGqAAvS4QpQUIk0pwnoCW2JyfbE2W0
niITS/+xxwpyaKBySbRn2l7I5VIgrDTnXAXwWy0G8nhN/YZtaGw7i6NrSHruk0L+EbmmZWDgcSVM
nLv8b20M4TvqhgH216KfQYDYJdgEAbfZggnbpvrzjT94TI81002UyiWCFkhK+XzsOTHt/z1ic+GA
qcdObobuwWe8y/qSi/z6RgjtCc0XxioIxwkrhiPfcSF5lqdrq1B6WyjLp3vTHM/78kJCLJZrDM2b
KikCA2KP28isSS3e4H9igsP+171d6c5XJ0EYeMRmlSw7Vibozp4+vJZR8UfGilS7S/MTmGIhHSXF
fG1JaOLY55TXNuFsQN94GydbSAabc9iKasGMRQ/754Qqy5aVflauJC2uD8SPQTSaJIdqwUF479Lv
AituEuex5ppfAnjYnOsW9zGlME/qe/XiSMYzDxitZPBknTPmQcja633XOLT/0xNLCMJteg/QDYk8
fanIS2F4ttJ2cVUlJeGxttuyJXak4ssxrSxrE3eyvjrNaUtJrykmq7xmYmamQjN7qKL9dVE4r/9O
Gh4f6HRp8yj27WVUNOMOGbX79bUWpe1gbUy08zDV6F4Z1fajYXRKRKdmZU5ftWF18K5ZqW11c3Ar
+JUcfZAruZngGK1Hk2roHvAIci1nyhceNvpNZKZSQqLRzAesUmXZbuFGJYrmEQzJ2MlrmsaqYT0M
VXQGqptGOuRijH1TkvOTqMSCaJblIQTNeOy3oqNjKAWFQPcuGuAUbqi9WznEpbZJ0OKAQKztPG43
rMTHTr8jpw5acP0HvekiuMm1ajfKf6QX4ef0aO+5Lw4i8DnmV7+ygeMJohRNnbKzPTXYTedlcBQM
kzkbKTAYd6iGSInp6X+c6Hfswgyyl0t/Zt+X1RqIc++wWRlcPnFPzujqZi882xs75Xyg376I9SZn
YVFvyybDyD6x3TUoyg2lBAqfYJB15/TkK6v0MDLRlwtBw8L4y1exDnZEFdis4EYIo/o72ScrIb67
vu4Q/JtH8Q4UumxeCEcYIfVDa05x22XRVfgGkqvQSB6SGFWwBf+LAfdYKIBhYRy7uvvwaDaJkUhp
W8wCrk4Kf7z813nwIWpaU4ljMKYUyb4f5sQkKlzg/xss0GL7TuTyakilEiVYnh1Spd5dul5ROtOv
gzEF5/m+Vu3TxZ3N21JYGzggAfy3O0YTOS63IE7gzeb0zEL4dv4/aAQaOOJOu3AUDQbX7aQomMt0
gihYsIKg47jmfXHJkENrOCaKVvw6iiXfqbSeV09Lb/LF4vDUMRK53o4fhfs4+v6RzdS0gxB5S5mF
g4xV2/oPteQsDTstEzVWE2B9xkZdBBed5U+pAXFJZRaorBksLxXKUQojr4Ry3CLpJhlA2SnlGgSm
1uehtSieaNpBHoH+i9MVEtTfkK1v0bRJsiTrAF6LA7gFNLMklNH9ICvR7FdVScdTrUcwtbkJCuID
kGwjRBQ5jtQXStYfkxoSQtdW0y1rwaMZvuehuCLN/oTLv/7qJWe6UEn2M1woUh4qECQbfE2srmh+
CzdaOysyQ0y1uf6MZZWz9jjRnDLPyb9Gt2QSUiee5+H2xMzm/6heJZ+doLxV00GT17GIP28wwpdW
HskZh8mMxPu0hdks2dx8/YjPeH7GMCLvsyh47LQ52R5phWJTliFoygIQmB9+657pOTyK38ZcvVHT
EiAMdJE4s7iHcxXpCQUMLf8wg9F/KXGiU6+0s9Rdpv8BimcuLetPbcPwGzhCJSBke5FgcVIRkdhs
tf4pwY8oN4ZXJ48/feEO0D/CkHg8pYJxLceq3nhrvnIjipOtQNs1JjElFdNmSTwmCkNyaZFqR6L2
rELMjEHizg541U3TCLoRW4aZ+qFpPzjZkGAOkmKb3FA2brDffPD/RE1836WiYW3cPQWFp4fbWK2d
aF2r6OO3zw/xLQ3wgmcuUlsh4BMB3zjI/eproCGEOmAp1LHawAyyxrBVvI7p34IItKqy+Nh4Ua5s
8YH4SNX9WAD5chRZ8UBy+GlrLZHhiixTFHOTpJxABIWsJNIFNaF7sy2c/I729Eag2pospc4vjhsQ
PLV6PchZgn1jTuALQG57qVIP8YWFjeqyr9XYfx4jvksm2bSVsLcdOU634I34ndQBoHMPzx2SGzY0
+OxxhTyDkgCuzHdwHVQbqwuTIXpctujxsF3hN0ZWdMW8d3Q8nU+TXOAnn+TLyYjJp0vMiIAIOIgr
io7VCYC2grcFn5+Lk82jQUtCkpJYfh8SH1b/vqiejIqgoFJKxaO9JRu+9MowH3dfIbP2NY1YItdB
K+ByE7XPN5YBer6M+z9NY3kXtt1uclCRh4PY+t7wBTsJqavj0fa4cY0DWIIcqmJ3cR4IWm1O3Xdt
1/C/faaZ0rYs9Ur2+x8OjrCmvpz1A2GzyVZc6g7gHOol2aEVy4nVsbbprtpK80gDFKY39+4sNMS5
JKC/ZRexBlMziQrE8ScNRujo3nBCJhFbUYQN5f5QzFSki/mYLvGfhmeEelqY/EtVFWlcZ6mKcTiy
EEEOPw2vmqU5ERSSmBZtPqxkStn+iXp9mpVyB3q23nvehKZhMDCms6I/2mEwsV14h3TOPd6cyd0T
3yM5wHQ71p8IyvZ2CxHdhnn6g8dF0OZP89Pl9Ao7aJQkEeiEe4d3F8lbD+HWjF9Q76fsOERfF45W
oAJKnp5KR1vnPxxsdh/DHKYCiFc0OjQiJui4sab8Ham0IZ4sfHoJO2nHmonxNyWgjV4KUNk6v++R
JGDXdi+g8uRASeVDn4xr9DM6BE16CuXFUJgbic81NvrG3xXilsWpuE8VTVr3v6d5n+2nI6FIG64i
eOfvWab7Hz8GdaS6/ATnsmrGCOwS722e4MKe0ed436D0PrTKUH/sL72LhY7jh82r+ewMXrgahHd1
nxHKFDdT7ZHw2tJlrVLHBdTiIAquJGdtVGGIAlZTa9nqFeLVgYvcVIttJ/B7gU5s/IMj6AGd4sbx
t/KZ6fEjgS43VG0UrmI8qwWNS5e5pFZffmzXJO4ZqWKBTbPglWDeFtjKmZEo/P7/M+kkH4yNDqbh
dp809PdCNGMciiJixxClIVzc2H8tpBIv1LFQZIL+14ZDsi3d0CAMpS0kP9nzSTEUfxZQ7D66+oNu
86HvCfckqQXS0R9W766zSseUKLymVW1hfdCU4vsX7wZ8ncgOfbaE5e8mc48tIRnNUpxIQa+M/Ymg
iD6GhhDzAGYcuHnkC28Awe2hhA0LPb4qQysUj1HFsSyzPZMo5OeDYQNDfKnobw73A55NG33hhNyy
AOxHnYL+mmQxKiHpTwgtWMleyAIvS4aOle+ILlDKyJTIdvuEnRCvGzpqxQM/21IXwUUZAWXaiF8u
RAJyvhZh3ViCTunfuk7IHTwFsJf6BOsX377B+EuXFemtISaSxGRX6MGOI5G/kLrRZ2ToBO/8/yjC
ahGY5chSb7Q9g5QLRdqaOrvlpuVT6c/7YMlGj1p0AlNMttFI4kejWsfBeHDsUYMNc0FnWGkixzSB
RCl1pclrHVnFEIgaZtn9CXHyhFIu7wqt1pCIsth2c1yLUemj9y+MDSn1md4srStnVM4b2Ye6p9oX
qwBxmAOIPCusx/xRlnNRixPc3U+zmZhs7tzWyN5zMsQprgVZVwKbwo5YFr/3nlJEOO0XcO20b6NW
xKya+N3iRpzI3mCJjlKYUTyjjDxDCJlZreZ6EC8meAIBOQCsX1vrYAOVe0Ab/X0QXOLOse/vX7NL
pl53IiQqMYbVCOl5hUbbo940SK4ezyr6YEA6fGR3g2iR/o9JAcXxuyOUlCKaAzTBeDC462WVJbpW
ZivG8wcRLBnhBmiwSac2xAhKSwpyiyPdSdWfZz53Pva/JYPgx+MwEeTXdVQY39ylcmymj7gxn2R7
nMmVv0k8CrdDryZ4u+bo45OUzgx8NnAqtwJZIATegM8MNPlvlldjz3R7pUM5I5k/wB1c9liSXgHi
CLMKQEtnV4bDy9sH/5qjjsR9JIllDGdGU84vz1pYadkF6YdKZG9ttJH7rXmTnfA/u+Eo2cl2RRsG
C5/5oNKd+Zyg6YesqYYKte+W1t7E09bex3+gixXG+ukfo34/CJnxa1WIg6RSdlcwrECqWezyfhyv
z5zmCxAY3sxr0I08M9V1ObFX8Q0iefN5Gyz3X3THj0OqAlYOKYAQQwnFkfhGUjgrFyWc0l0i6yLy
5NzLNgr4WqPPUTvC6K+yYWNZsdm77GiL7yNKpKwoLBfOMaonYj4QJeURSh01cp4jD8L50q+Xkw0l
2k+jWCQXdrXT9xhYfj2uQtDvj+zfI5tdpqkhs9E+u32tlJLR0UTNhvphq4+7RrNs83bpMgTGQmF1
uzStkQVdSECvEnr8d29LM5XDtplf0zIqd6T24vUl6Z4NutDVTFRvykuueulP/1AwfGEohV3bCBal
+cuM3YUJc84KPX/3pJGvTwmEI7igk2jIQJZMbyfN0eNxWTNUwpE7ZriFDY4LG8c5IM6FbGFvqFA6
GFb8NWqIdo+WtJ0hhmTfJ0HAZDW957zDTZI8KUjf0sUrM5fa44CBUamF1tfeVg5xsSY3riRUVBZR
0yCY+z5z3dFv8wUviMToYwKNOzHI/SfdreSmj8zXGPShjr4LdHs6t72BNYjThRabhwcXFFswP/dJ
IsDUxwqWBB8jVxpGIFH2j6bqgmFOwc2qKaeNJ78FZbQRcl6XWUTN7PM8nioe6wU89743ijuJjeqM
zhH3fSEyaAo/XzTQ7D3Wd5tXnnsqmn7og3EDAZ2ED97ooD4fgYzXZzmrZll8VPOLYFGcFhBk4S38
834maItWZc/dLRQXnKBT3MkqMfTqMquq2XMklxHJmfFreeUVyHlccByhCN7SVthz7P9bEKCMme03
5s+9hCDLVEyLXKwsQhO9PJ7q0ljArG5RKukguAar2wQ5myquMmEzWHB+bSidwnEMr69lmIDg9lZM
DXCVOjjDT602WROg2q97V8mz4XpyrCZ+ViIQlL30l0SkpDnDMbiDPLaNcRRd9g6cVk1A6hn6OQLS
sLFtBO5xC7RdYzFvXtYXfor2vkAA/8zouIZDJSzcj/KesT8Cn4Tco6DVBa1sY0DmbRr0K9UXjdOI
/DOE1or3HWCm7YgitgByXXBvOPR5kid0MZr6Nw//5mOkbOkUi5Nnl5l5I0SKXGZt4ksSP9a53QN6
yh2reQQqIVGxOGIYLuIiMAPz7TtjsTc4iAB3m9hH0rnHie1XqvdfM48p+pM7xYBAoz7Auc/oibDW
vFn+zViYmSjt/d96NHzOwKn82eLV7DZLEq+HeCx8GO2qwkSaRrno5Li6wMCip0fqscXTWDJPK02Y
ca8G4OuUoGetNNovZ4H7JN9gh6itxXkylmwXMUO18r4DihxXuiOYuOqTJ3CVBy3LOUl4Pv9wABD/
KujzUiHbm0BRdVgzZAgiKzvRZ6LbgcWUR1YTPXdI2/+Y5TBj9EM8yJe5j+ifTWgEqwyNgigEFT7m
Sn5ipIFmbId6B4NcsNV7weMhtWNUV+0wIpfvNBTwOiU/sXzuDjMHqfITSLFZIa+lxPP8UEcpro8Q
M8qjt7nl8t823w7w6xAqZdP1xSjZyAnP2ihiw7NJ+ojsJ7r7BJQbM6biIZnPit5iTahj9lQ+QncX
+HzQW+kakdoLqhDZPXYMN2CBR362Fz2crD5aIdBkSTPZr5Bk8B4uBF2LAzuedlh2+zWIZkWJdUCP
pzptmWjOJcQdWhJ9XyTl1ZgOGJmB56rNIJ3v8i7DxlluIvcPMLH3VMZcluaWxwXzpTdVUt9YJ9Nr
6PWkih/j50izG9hnc0lpMfhcjXWEz/AruIG7XdFMBG0WdJW6nqu+eldUcDK4A18vaWk7PZUPPPK9
v8yh7GDQZ+adetWf9yulapPDYhyvuaCczkMKr/2ktOMzS1ntVIhgKNba0ClwSn9pHPYXul+FHdnW
D/aGku+gBssxD8i3RwpcTGflYw1O3qI8FbKHBv6uQaU3E0oWs5YuHFiA2JmNsEZrWNtqkvcDJDSj
2cg5JeeEL+NhwdsG8i7hVFvQQ6IXWzraftWzsSXDauEq7VRGipvbB7i+hcYv5gCwa2/k4TxF9Y4c
XtbVjVL3+tVSZxWRugQ0H9q6MnKZYyx/dWYg0DlCj6yiWqGbFoBNh5+JaLp76VYBPeuwfM2+lbvg
DkpvvWBvrOLzrk/llFN2n6rGVSdYQHi1b3YlKgqYbC4GejrfgtgjDM81VNf1BihHPuj7+k2HCgSF
+mfgYbWgba5pG5yDfm/B512WpQy0Wu7BnXJLAV+DKFnxEEP5DnCIv7NP9ZGVjuvx3LfPDbEv/Aj0
pkBy+ijlKQu32HLh+87JSrCruxeykywgrrbEMap6vx0h+9KIZXP6GZGim5mNLfW05erGgl2/nxtb
UrBbLKOa3kemqrq6RZ/w8qKKhOfrjPbMJigNS5On/NvtDmSEyE2q3tcxTUAtlFoJjflb9qJ3cAIj
1R5IOqLW/m2V2MydxSPdJGGrXim3pu7VnbaEUqk+Yth4GCZz8uuqJgggmJhCuzYluvec6V64baf9
nBS1z2IE8ZgdeJRL12FIRnoHTFPCPZumZ2r2/fiSrwwH/Dn1Y+q+V04oBqL9aRiwQr7dPdB/FgzS
FUdHkYuSyY9ArZwRft+mH7Ek4PZwuGZ1VN1IiLEQlTkLb6Gs60LeljQOWOrorb/ktwsrKtbN2h9r
NnYjv/NFjDmAxUZkmBmfKXkzFioHxgxLCkgR6mc4UZlCfxm8Y1iH5E402r/138U+FHtOEyAxoRQ/
wudcWKReeDnm8e1IeY6YQN4T4mdoCBSZn58oR2kAcIZoW9GuJYyLy76eseDLhA3CAgF+0eNKnwzE
lSeaBoClXwqddpkqOA+hmyzu/0jn6oVl+0oz/A6xENH35kTUEhR0grsceLk3EZ+2sXGAya76+BGa
MAo1YvzHmQkp9S2Xlq9Ke4SqqEtKhYlmRbC+gJHL/NPsubznS7XZQtmV/CUY+huShmr0+nlEnS7n
m2IqpNqGQUIYNl8ebx179cGwggYu1ON/II2HAqZQJCGPFmmyb4SQfG8l+6Nss6bM72pgyf5o9POD
LX6R8cKBkc8aa9BgE413ZpTxJtpJ0H9fU0VDizNnUsZcAaF37mwfm/V3/S5t7kmWVETuwl4pu7JB
WEzxCjMQf52xZxWZ0u3EmjMgo5Acf/ENTTlHos8MEWLW1A98KgmUn7Twhmz5pTuD8vRXEbOCXVLz
XkM3ukYDuh/O3wE46AyuqESWbTqn1cTzoatink2OszH0MiBGrxt1KmoVZg8RnLzK5Q2D7ryxw3xT
hgj51sBl/lMnVDGYdnxlYr9ttpduvoJcwbPDMEbmOSSPaqSHctuuAt3430qK5LYqKvMhFH2DtaFx
hpGMcZb1/ewojNfCVvUJjpcYKGVxTXzn9pn+qC+s9AVRUHzbx34N9sN2GTL0DFoPMdJ+CJ9Oi3Iw
P4dP1qcZH1Utg5hMFheV0CtxbATXInZ49z6omcYDaCkqerIwsmAoFYAUAZt66ilq9C6wArZSl7h7
9LgTUHpkw1MFOyDC04QzVlZMa6tyR3uIrJhzZDQFFjXAV4FWBYVsL8LdNSdOeGOntM4vr3TM9Nke
x/9UJlh1YU7DPOmnt3+092SST8o3xXMFLRBZcFWvMcag+UjGfmWl07/MgvHAf3y3Qi8pSMLsxYiy
k4oQW2d8IcFJLCQrxXnLdldtBeFgPYKiJLeWKy3p9Er2Zr3BdCNzW29nTLAtj/FRlskbEUt3U1bZ
pAIqeI2Onb+5TAQ1yn4b1b5o0gEeI/GbFmzS8NbCXv9IxVrnh7n93JSL5PW04EeaOfvs9H+FYpRx
J6U+DiaoU0+TQ4GBcLHOTziyPPxzybQajkCc2XG/GLhw0RCpz2ZpWi/LSrPdBXsUbEeVlDBm05ow
oEnv8e1TjVcdi4EozIaXEkIuiR+GQvR6y78FYAS3Gv/JZ9mAcW5yXuVL8MNUUqEdBbatl+bAzKtj
9AsnTF/74ubg4bNX2ECHRVf01YaR6YtjpfqEeAOdzx+NhrZkW9j+IFMbfn4I5eChAAlGgmq5DfEt
e3h/12qTWtZCs1q0o1CDdkxsUaYpF5EJ24QgjPkaJZ3YNnUkNn8IuI3u0G2JDxRXfKkc4DEp7RgV
9gzTwXdSWQn/+LOr2jZ9uxKQGyOtx1h95JaEOXdY9EwbBWXCI2uUvRkaG5DpBDvL9PuEmIzewrcg
kwhYZrYBx+qMNMcWWlnjc0vs+2LI5faOWXuaqcgKVXNvqU0GYq6KiXGSanzfDKcd+bua4m6/USSv
hIrlOg7n6IziqgV7RiHL3hX+/dihHULP/SMlwMjErcS1UqixNGjp0M/JHk83s3j7nLrYyZDgE2rK
VnZpZBA5KCkMBsQkX+x9/nLUWrRHLWnz5ZbgmTDgYX+ARqN/d2MVAUCMhQVGGupEEafs8fBDAAIv
WgyFB2R2jZRSF4bFJVY8Z3RfhNoY5BlVsWYUDXFRFp5eSRULqAIUOBEP6xlqddnaHekCEZYvNM3O
kfYb3cR2xCfvleseADCBIeVcW19AyJGKb0RfJIpt/FtWwLZeh9ZbxfkyP5mX3G0G+xmBa+UkYe7q
S9z64q6akR4/aK2wY49fCKqxghl3giapb3lrpwDzLMvnDDZwQlyUwV/Kpus8ZzPnu+tl14KT3+ib
qbSg6UX4lHQX+NM6x20baqKzj/TafEN/YWloNiM49w52prtvf9e06qLZvD2x19uy9dXPGRytIucn
RMa/FYMj7V0+7JnwtHhE2E7o8VljftUy1V9OBdSLW4OtvnfcUY+X0qJTuWPeaN0Zg5AG80RNFiXJ
vhOXR2xXcl+csoyYoE3e1si+VxmfWeY0kKStGRifykNsCMzBRVKXIAP2C0RMoci91Zv8rGD+Iyco
eh9/d4P077lI8h+uDitniqZtlz7Yv4xNloeTMuCr/76gCRiHNl0/g3KQ1P/iJ19rCdMtKX1FnyOr
Rr8A2bYJVXxLj0z7x6EKi0GmjqisXtrc9T4+qZDUYzCgkyGaDcbt9SQL3W2hWVKpupQ+p7JkZ6pD
l9e8eiUuTHvYUOekB/mFPsmcIoQMw8pg0uxLdnK00ttauDNprsT/0d7/Xqyk7m93um49OK85M4D0
gUs72pzqE/nP8VWiPaOVpDnuMUUkNbQ7lw8eLlEfDUBxMo1IaYtaRIWki7q5t+B1CmcPEw8ocM5a
jEJ2uEqISCl4v6iXKkwuUdsjcNblxml44Aav2OQaJAhWbzvhstNGOC6B0K7QZ1/f/NNCADgCV1po
u0VgbPUX9dC9NqOJX6ELN/6ALYtQn1d/huWAbOiLqRuvE0qav//ZKPAqeNpRzhvQs/F1YX642A9V
Vlw/XKVEjENsrRwXFt5fEcnyT5bsOEJcEmwfD9Y/dZMdldC9p5y0g/jJW9kf1A55/ABtTaPkPuWy
vD+QERDG0SaLZvL3D6mYMFrrJ4vkzoQ4Gv7L4FpalSIRxpCaVdVUry7E8EWKSYeHv92XWfBYxhsA
3IqsQb2KVau42fgsNmpkBj3DelfLEY5AJPIM3e/LMu+1d+kBRXLGr8arhRNuBaFj/J+vanJu0kSR
2AhdkL3//738iY97IchSPcedh76g/I24tCXhqDPA9tDUyJSgFcUTYobV/o5QfMupC/ECUBGPqsVn
lp70r6zJwF981ICtiqkMPj3OfCYeXcZq4NyGK1T/ssGh9WfNwo/7zg8Xa/GjTHM1Zf7rDRDH5Jmx
/gdUzxYxOoW1jAFNSoky1+GE2VXQ+uqThgtNVO3QKDnV9TrhLMQWiJEuVMBlAYf+i4i5yOdJYQmn
j1lmx8FjCJDcCJyEQucq1noppFZzJJYyXaM4x6UX9ButwfFawzHLfM+zTx8M7FNiVcJDeYGZCQVz
WuGfffckkZxBtligX9IeDM2M2N2XcbXBIzRYbP0+fUbcZGcQolBDqfZWFCH8BRo6j5I1BjXazYC6
XAjbtOQ0l2FZWKRzP75Um/sA4liopPu2dBgO/SNRYlc9FZw/3RpavS9UlSnDOqXhs+Qufeeh5Dim
hMX8hBJCvD+GeT8KKlWHBbixLDc5QTrTxoHX0go3Hyj0lXGoLkTi3VTwlN6WKAlirHucy9aa6IRw
Z5x51eI3GOV2nEyRjqQ3DsMxSU2Au47xyFTuSkAQ57UWK8sQNFYFbv/P0IRhNPELd00wcxGF6URI
SAlwgvY3C2z3LdM/kLAe6wyrQ+j0Fxwm9ATNmWO65E8BpgzmSJrsZmMZE+GmbFdC0fx0M21bRSMT
g7RzRM3kJ0cTa72V4ePilCKAY50klrl4OfMpb6MiN3dYldMpCIKXTZu5JWEuD98dsVqbB9n3fzln
zjA11Hor5AWaFj9oiKOiVzdooS2C0av3cqMFEwGrxuNx469JNZ8cnGYNaalXwTCmonlSP9/3/Gwr
TdxF35fl/Wx2ZKaNxpnDcGlQUN40GeErrL9j+dgPenmHYZAtWkvIHv5xGTxM1J6eATRciSuA7tQe
D9WLIbVVzV2MW43ZnviUyf0szZNQgI8Ua4zWKIPyXJCFg+CYGitUJEXf06NQF5u+r651isv8Gl9m
DemY3PhGgUjCMkAlxg+DTgcNfZnbK8U+A/L86ywDOIib2XZoCwSn68dtanyBF12LjvkQtSA4U96M
MxrvFNSg6z97Ub2+kTbGifPR9cnzJszcFJDuW0bwwHOHRr/vDFEb0dZIwZKVzPhctOAXe5DBlA1X
0ycAL7c59ksl7mtrFHngSuPLzRI+jhV/t8QZbWSZPj47jMuzb5ipIjDSCGHaPZg1SM4yMmhfmBo3
jUMB93p9CwZzKmLew/z0UhBsx7v+nyxaKrAlUAbn0wia1R8OL9IX4GNVhdKrUw6CV/O4xQlE3pfG
6/dWVpG7rSBYUTY9MUCLQUfiI8SOQm4GS51zwMjYMIgPKql/wOONS/GNtFEkVfNx60Fk01L20cfR
+0hMBaAW6qrZiSIgfF35fWNOUpoIV1Nza1f0uc34LNlAD6Sy1lyCryyhWA9WRLBaAhgmmRCPU8lk
yhmDGM7qmFfQah4xPb+O/EzyVU4IVMW+SdKCq9kw0WPzBTvjGe2k97pjtVzUqAy/C8LuRwF9sD3l
4jOCFV7oX67X1e0YDMSJQicxilmZ9hhI2Pxqwif9H9zdelqaJOKMb65XCunSS9XF42v9Kgyt4uYJ
4GtZoq8+37xFsljbBvOL6KeKxMlBXQPpusIo1C2F6D/Cv2/LmJfqZoJ1AxFMl3d3OtvktCzIeqRZ
2iUBMx4vUL1JLee3BTyWdNlJyn4MBn26rJ/2zts4S2C6e63sUNO7APjA5LbqWHxnsaF6ywrpII9o
8ZrjfHh/sAa7SbiPdo6pIShFKnHf99u4u7T+m9mYffg2rNZwNlNBuH3iHOqiRxL/kaocrhcQyAaA
YQZjNAepieA/1Ww96nnSR7pNShnIm8T2Rt5/KiVw6HnRnaL34D/XEWI4zi3Dyd/B2T/CwdaQaLWG
/KJBvKZjkdegvpn4u2LI7g7PZzKEQ9U9OozZjgrmQinaKN4WUF2CPU2LiTdBVW24QiZMmcCqb9ug
Eag7R6boAO9pxtKBG5ejpPaHy1IYK3vvUGrfsLXCoFGS9pkzJctoH5ig/SRzmofrOQRxZqaUvoVv
ygsh+SR0Kf4IZEpb/n0nPJoPXGJDDfJVgK+en/mpZSJmtm/8dmnr2rrcayIHnEXFx2+74dFJNPwd
veml7rL3sTCGcCzGojSdgZ/as1ghAlVIDA/0LL/SRq3PW4GUtRStqVxdQLgkgNvI324yZpGRTcpk
x8L46ohJLMoYvCQHkvG003QhRjXgnbjPnsz36vRmBE95hBia0kzcH/s25OllnjGxhUfgaR5aab89
BIe1SfgKnXvMC1ucjklUf5tRAmWeqsEIdmOVwtmp89Ma0u7zhV/4m06jQ12wUN4QC1XgNTF+bQp4
3jhNQhkZcQKYCSMEtpRu3/4ELSVR9VVAdKrYtCqSp5ZcZuW4sUQPB+vnwtaNJIM/Sqkx8BmNXESV
7MSK06MHYoXXw0HFKdl8YYLaeYl7JcN31XRGJ9thrNTGBWzsFD+n4TgjFm69Iioiq1grCXW8S9+i
bhOSntADcTgxVMXUMPX3350t7OMEowwreMH0g8yr7Ig0gDCEEjk5NwuWnZl2dcw6EVGyKJS4PP/1
TToA43+7DKCGUjOCUQZw2mNMlFBnJpnG7uP19FR7dIrl65ITTMpH3RP/VTdsrU1VaaAEe/OyIOMd
mFvbnueMAHbR5P5TPuZAw8RwzqXOfWTry1aBjGYacJicml1LYr3Pzjfnn2aGxAQxgAYqC8/ThL3K
X0nMRvbDI5f5HCRptyDoqty7DpDxg/gtd3DAeogy/PX6V5nSax4WkWY3CG8+PWu3UoRXWXS6SyV+
hHdUdFO4NG+dE74H4Ao1huk+wx61tsyRot1GMrl1E3qQ6jWqkHW8cV/e3D/Nvpj/rgcEzNTQ/gaU
g1zv2zukZsZtc/DIPeTRAPrq1mWWsFBcKLiJM9qaHXWihWDtXGKD2n9eUE2GxYJkpqTwN5m5FLSc
tovCfSlrgQZU58EMdMufl0Q//1npHAeN/aEZDyreOKntoUXY6eaEn8h47ouIzavMq3HDtJrS/7qX
pIFpi7fUcUlr/tPO/sXQOf+Wmh5S3Ja57NbxCxM8Ce16F2xoczsBODP/KlZWIoDObU6FcCIm/ufI
W1X2UypO4qWr7Qml1jFXvQH4NpkTXFJmyQXE5vGEW7PkpC1YjJKm8zpI9Mj7YiHulX8oDoQnIpiS
0mYwyarz9XBbv/Ql0PasdOfaq6OVBByr5RXlHRTWjmWnR6Np6P8MfSQNq7fsaFXvRCDa5fXecYG2
cghTT1mah4IekqfKOO34n/4OVzWDyGuqb3vfLrRHCRaE9jTPyuD8TPUEy1HKVyn3BLCuoOx37B6u
di0F3BKFUMdglHowown4rtmi9YCtk/0rYNkPMkAlgawyLNzS5oGV2UrzML4JJqVeI5cDo/m9cWsM
/vfDPivjavpy2JL9nJp2qjt2pND6IdvmpAwgBeQ/GZAffu4FTcy2a4hjOojxWdOWoeFikLgu1e03
qtMSYusb8xJqumeSEsOb6zFmlcs0W+ePLX0+oCOovL6OQtC+EWjgSFq39cqSW3rLSHb8ZPsluW2h
xKReZi3KwT/ICjQ/avV1DgoBcAdEavnjWhj/yYtNY9NNFJD7ZMZiGGejHCYjUw6fbLXGL1THoMeL
tqjK7X1TAL81t3qxsVP3wQI4niFWrmAiN3cAEQxJcDlSSaBtgG3hBPhc+BJGVHDXhunhLALqNPuT
HKGV0vrf/64qUp59rdkipMbg4vaF5YABVnqFZ5zIL+ApkXGvyILmMPw5mI/JeUtUNgShd5TLloZs
S4AS5OfKb5EcNT/wzpHMWF/UJphJzDwngIphTVoFkiCpLpqMhtjl8z7umWPp9dhTQOkKp9vRApLw
4QfDNL4r7Qwdo8+PxwbqC8dp5zvUpu/CXk+dSZV0se1Mnv9ZD+UFFZ38nO4q2UhB6nEWoT8+h1HB
wK8X3s5CeZFF3lbhtb2+5j03tsw6YnPpHBkdN6qifdM5EAgS2/3yN86STRNpQF//1nG1c4zwQndv
Qgrni3yKCk2UU6pj/Zm1MAk6R1poKYGBvFJr9jWHXgEU05tBW64BodnQ8bodjPm/LdtLA40DyYwe
OA0f1lH4YrQE5XxGXz+iw/qPGY9tpgeSEFPlbFKiyzzjX029GfWO9MvNo+PnPw0qrQflFgUGMeVw
FcoV8ZM6vPwTE7yqvU3gpcxZtYmxTlP3Rk6AeOHaI+tXof6VIqy8L5LxBLgXeuJWVIKI++vlQZpo
EP+2cqI8gqvpRj85ggbUfBJVqj8oU1E/fcWeTeIm96iKgasHK7CQZxlnB7vjaF1MbqMnePx+TNWC
XETeTiIaNK/xjgoTBGkJn5AVVWA5YEuYOWq1x+g0XNvimuxklgtJFytZTPAcXb9K59Y2yDtv4nzr
mZRgzl/jkgZIoo7on73tYee9nUbM8RzNrYJIFJ7YEVz0wnjsLrwqGyZxZkWYSSfutO+JN144OJvh
YLgWwJn0iNgETa6niUtbqtqroUrCzzRl6RbT8SSDR8AMj4ox1bG95A3zS3SoDZOxhWr4/Md2qEUj
Z2UITtNrps6+SOEZC8JYrybhqX22DnMpo489LSiX0q17UVG6lBEf0bUvY7gg7lRcYIGU1Svl/wjO
4aSkh9kJLSJxHswYa6ek/mDHc7cOSHiF0yiWm46w7dOKi0EbD6KRZZzh2p3Ntn/ez4RBVA3uLNLb
Aswq673pAGklhdS5e3597CbzGbCfk4HkBLwyJp+S5xCqYM3YM+nuykBn4It1oCaLEqMWK6M03sOr
E5DtE/u1w2Nb3l5M6dtOB5caOwvRpUfW378ZCbF1O6TA5tWfRnPWdCEZf9XpiVb1hYoBqfaOYq1j
s6RUHKvc14XwPGP1V5xo1scKIp7AQ9PEGlEGa9/CtkIC+ddQR2oh3zRsirrcAqIlgcq8Eb1hNSeJ
WbOzSQVvAfPqi0YEDQ9RCYgUkp88X1aMeVIMYYd/bC35kL3vKWJpW4pvpaJ3wPN6SfjLjyqi602O
p2kAxadDsYkBxUezBDrMkx7h4cNwfY/kfIXfukS9biUVkKwVPNpS8nAQysiKYlTp/5AkKCjUutJ8
Yqps9VGc+clKZVzyVZaXcKq2k04mRieTZQs4ejwb+Fw1HS02lJn3BtU/PDqGtmNyjnNIvHQ0Qx5+
QtshHewSW7a4jfn5A1LAficDmMXCcWZHx18BWfyr0nK8LZ2eJgEZiIuRO8x4Mfw8q8LnbRZmVj29
LkSB+QCKYUPmrhqigg16prhdMZDuNAUeRa1asrTCNP3YQ9iF04/hlEgoZPn9YHLGO/JexBhslfuI
IAbQhVOh46I73rvA3nmIeBXXGqRnMyLaWbvTEvw+eyFz6ezFKi8Eh2jD3uGUGM9PBMIkt4uw//Bq
3DqiwhwrMt594QKQC8RjNcbzDdFT3pbM3lDOGjsIHilpxdZMoMpgqiUJusW7v76EZIjLsZZNddbT
BQEKu3rer18x2ZQcaXWwMn8FZUMHn5fmwHpofp/FT5EUPpNOltXkOjrSyX2/uxCNhOH6azBOi7tD
+Br4LaSzpEAo5kErQMEQx1Jqi1ib6HuGVeJa4jrG34REWy/21wlM97zI6PcBbxgRVqGo5KBuu7EI
7gQe4QPmmmNzsdbQEgVsDsY3v0nWF1CewMHs23uCPkrPQ1iQQ3hqFjn61e1A+WG6ZcQm0cGm6e79
zZ3T1YEtMc21rO9Y5FbomxC2JjTElErxzp8M5q/qk4JKF5yrtxuPFzewhLjRS/i9pSgpTntweoPn
huQkzehUrZfk6+ax0IsA0gWiZ86Phees2K9FyHqU6XRqgQeB1hE3y9DCY1+tLFGWh510TFhPibUe
5j/outryni8//VJLMuaRBy/m8Gu2eTnE6XZLQpSkkJUqczHPH/7cGrzn2zRQBz9kFiSpH5Km4bFR
NzQ12JwY054nvhOIA16c0FSOX5OkWjD60tJuNPUpjn5RFlL+pryNdkAjbFxxmJMRARAQiSs3vvKQ
zT9tILrnfUguwgUH+PbSpzX70n74jlGk8sZWt7rn3PD4SUVCd0bc9gDZ61eREYa+rDyvqZ4MJHNs
v/tn5WAAc7jCW7I53JjDTBl2rXqrqQOAWSB30v7ddtz37mfGcxbTE688kf3RYO+LIWi2rZQ8Hq4X
FyYfQXRhqNcSYfGL9nVkE3tlWe7H2r0ajITl3dULOXR5ATI26NhfwCcrrPeCGQ1v0m5vDKTvt1Qp
IjyA9w5Hzp27qTJqYLtXgDDDbAuTzo2y0MdFi4gY83YtA+jqDcXITbUbg2wH6X7ZCYHqJNbmxFD7
yVnLOwhvQp3L9AUJOWXMAkw/eYm+9939XWNW7PNuQ8rDIH/emsx8zmAoDoo7JfW5oNK74v9b6RvD
4ngyR+Sh28q9loKmDzn80Ll5er0dgIUj7Y+PU1+ao1MCayI7PG6GdJOqhPYBEBRnBPLse6CxzuBM
NYGso8MBICmcEXqIDy/e55Zt27X+tRoQ4OvfCqvATi5at2bcPdaLwS2A37wghty9esYy7G5pyFw2
qd3JXVm/sXzRo8laE3cWfJe9/P+gWHL14Eui0PLafKzMqgCaMTmcoucvy9XToMWOTpn4HoES3yYj
gjU/TtjGA2cn2KP2ZsXu/Cdxxz/xHqsQSD6ASqUmrevd1JTt5ehcru4hVY3ir2navJo4Dg4cgN1P
M59hLrADNOwgSd4uoC1q+TgZDrFPMW3d66OA8XmpI5XWeCYOp66AyksLYjYI/3EQC0v7YQRqoMsn
n+jdP4vWaVciJrFiUy4m6q7OLiSq5Kd+UruBToq/UUk8y1xkeSFUANWdSNs6OENl5jETekpaov9P
WqcFM/nrPrLTrtCl0zks4l8Y4n5IJ/kinXPcNShwui6rf85sA3A6FXvrvi9iusDmFzjGh0AB0Dp7
aqgYCF/vCMByJu7drjBCf9x/wxnigdtNFf0VFfyKfXCSA1ekOHm9sMe18jGSkOU+LNkExCsvylo3
Y3PSGQzjkv1RHE0HA1rUTWEpV9Rj9tfto8lb9gt3iaiLgIWpVBPJ4AS17Rd2PoHCjPjDskMANXid
LgSeMMoPjq7VqzJpG2UZg/58/F55VXhNE0UuJkik86CjhK6WS5ddSVH0Kbq0iz2hpBUVrGQIX+He
7RcI4d7SuqFRnJAdKHqhqpgMBAZVJ4W4mvJdaXlqiCe7VS9sEQOkHTCcIhgbuVz3uTj+dDa665LU
mPnUlkKsZMaYWAjdPswJFag9NkWNpKzIAmN+Fp+tW/Okc/+JaSzV6N9KUzaZtrV75ZLgk8WL38qD
1OX/ZdP7VvGjw6DcgbUEWDdACoIPaM/IbIt0RbejJGlOruCTM/fm7J7bNidBkWp6jxOpjiQCcwAL
ZkxbjC/9f5PSG0U3Ls9idb5a8TxYW9LOFL4n3UJ8z9W2OMiy13wLtEBCcMCDSpLb2pu3mQQLhisz
zhtmgWsS82s3lmBKEH1Yj0Qn00bAhy4bJpqU3xKHZr/Upuv45x6HvZC9APfBZUSAAv9NjagADIV5
Ukgsn20UmFB5HEV6Z8AW1lsEbcHeMFFdCS0r7tSxK0R1r2npe+aM8CpT3vjAnDKAsFr6xG3lI1fo
IRpnvfWxRFY/svndoVzQ6EBHC66tfy3t/7OjVsprg4GEj1tqoEzdHgfajI/xGkwzBj8Oq9O/8Izv
mwldSK6/YyKlrXTMIZEgsetTIC+uW6Smg8NKDKXg7DlwB3PmmuzxJ9q1Zm2mQlVU3ia1EhRkkMZ6
B/93g2H7shKgaeZTaExPCbQXxrHgec8xwaOaJOCA5DBreACBrDppNcVrM5BaXyLfipXQi6EMA81I
QTDplU68+RdZ5hRAsBfKPsijOcx6xK9pIOqhwSVHmGZ46pdsXX00Y5HUTGdhRNkCaL9DzSr74QSR
f+iWol7ekDVB9KQ6Hf1JFdfxYwBavXmfn3l0lEe1gKKcIszptgiPJBg5QO3lWETeWf3Ld34aLfJ6
cGsP9F3SB7e3h2CA6Pl7umOFI861xJOaWvnzKX7L2Yqoh38d8YwBX1N+wBi++PJCwUS/4nNnK41Z
vlhs/+odMv00cmnYNPXjAjpTkINeJcLtG8sHl9DDUDEv1J/fYwqzdJslDflW7LQ2YMaDFtJN91Hl
ZzRA8Btgzjfkg1qEIVYwzEDd++8rA6UKimu4X/epnn1NsKNdy1Bo+513UR+DaAQgGgsyntwOslZ2
2K5gBotgh243E9TcDfbItxzzKK1FfZZIXVqx/T5iKTRuTLT6fGiK9/WRzuGhkDeZb5vkrcK0OFzS
BCrnrNJ2rjVT5Aomx6RVqccRu+OS/wgt+JyA/XD4W6pKQKmQs4H2Mg//EOOaEdCP1J161SWGxJW1
OmpgGn1eFfBVYNyX7PjCPf+JPqHQIz06Aidae9JM3lxIvzMrgm/WfdKWkydvZpUvVNi+R2bBDAkc
s2VUPpiv2g0ywWujyDkW/oJ5i1DGKIK3NiA5mP9ODuZAe41kIeMlaSD1DiKRm6++rfP3sYSUWWYx
BUvpCOMKvgCaen/5/jLHRHBX2ClU2JaCFn8fp4WqY0OuyHkUq9JqtPxU5iCAqgJcVv0Sz5005AyZ
iVFSxpSFPCv6PL8/AhytvLStTBDeSTtNc+SinnG3b838LqW5KsCtfyWhx66fAvIOu4lhM9JsLTIa
lx0rBEQsQHhWv637JA5dpuv//hIojJpWzjTans0AvxXf1u869VleU+VsqOeXKkXI0TN5j2Z7mjfr
Bl0b0+K1G4HevL8sluq1P/TyFo/zw62ohIlF5JBIjPqvWlco9Pfrt+Lv876t/sAe+2w/S9QStz3g
ojWAWmwSnnBYQ7xDBMIEw0EBTtAntupX5muNPRdT3bMj9eesZSC9PWsaccsYmA1sfihDHkrWShNC
w3Arf1Nf7f8pph5sXkaO4vUZjkThrSpnlfRd8vt492UvaVwLspWrCmDRNVTMbJRZVd4VVWRnbK2Z
D5kF9EqfegHJ28NeSC1CzX/Hf19iDIT1HuAqUgoOOa9vrPTG7sACbTNxIpfeQrvLDdqOtEx1gVy/
/yLyyom8vLNdZCa73hKiRXP1C9QJVBvw6E735R8MuhfZKE2PwbTqqowQr8skRUWdNqRgAoJPbOYH
XOZ9fz3O4Z0DcBNDDa3WhZc0mGb1C8OfiN4yXl6KArH275XFDKzzleICNnphgj/CuoYwtTelnhI5
buCodcG+mY0l5wPymtHJEXQknqcFLl3mqJDxkFyG2LmGKFp+fzMiTJSWeiJRX2sqRF7tDwCG02fR
YrTpcuhpz2piCUvDMVZ5D8a//j2B+ezQ0soFMo4anbovsKUpuSjLULbaNBK5fig2N9impVlRJN4y
lthZz1ZWEVCRkSW/YfjvYFTRUmiXud0t+KJmAmOrcjsgUwGOYzDcCln9c3UjUxFdek8IaX426oQC
hXDnFa/CA3mATCoXICjYYqs1lglhfJOiryu9A/efTjgSYNfSakzyfEJKZCTWmSQKTuYOzj672eVb
ZcuZXu6v3l92RdvuYeIpaavHfK3jFAaVkOONac03jbcQ4hCpkRQXTnaXNd1RLeBnQzutbdbjI0Ip
OHE4I/twHsLXCVo4/1VzsjAttSQkTAAn8gKPfbdAtrCNTRkfhw5I+lO+058bVK9Be11xNdDdVX+6
hl4LffMn+p48vcF3dto7oIgbhAgWgG2uphmLcK4Rj4HwKyJpDBijvyUUEI9SANJZaUxklcgS98CE
ty8qf0NfLuLvNu8VHLcl3+zvYW7KM8/UufUDHgNCGCrZ0Ugb2yEgG2ZheDn3bvraxPsT67OWPnyl
HlTaC5JNdUBStCjDVb1MqE2cHfXj8XrEECQin/YKiDsySofIi5ZHEX9eW7yBKq6/EOgLoiK2fqWN
LdXQR6fKuAyVbX654gBwXOjViviOCZeV2K2hIGxaHbEJihOYz2ZNEf9ovJF19Nva88zmNltb5raV
wxIWx0t/Ye5ZJBQazTeHyZeFMBQjoJxi08bAkVG7qYa3+NpEfF1dHmjX6/M+//QWT5Qs/UZtnzw5
FcQTsbXgFlGOwFEHcwOljnk5pW0dbR9K81A0LVQMfJ/qQspbwZlCTcnhERk6BkJzM/syEqsAVwBw
LiK2Hda9erOJ002OjWtvqrO9jNhJ3n+c5fuQn6Sz7Mub6yDvBXJEz9COd5kDFPL0uQG8taGyJ/Ul
e+rP4E9C1N1MzbZ/9u55W7zTWn4mB39Z8uf+YVcXw6AefqtANIZ8KN+jTZoTOAok/nFuR/HP1NkD
G9+ntgA1lTh48gh7sPUIDhfA8IKS5LPBjaC79zDQP6iae58w3ZWiptwj91qGyXFWFEDeomNQyhJO
e3i6wp4SLkfJawgGKcizAEWX0X/QDacxFw/sZH3OivUYDeMqsvP0k3Qs3rjGg90xdHxeKVDACdor
MCWTvmRNPhFGpjX3p0K2+L1qSaT31m7Kv6GiYGkCyBUg67NOuTehc9cp6nq5jWVjOQXZzLSWzu9O
YaBivSTkWRzdzR+20cuLUmq0V3rvRWQWjuh2fPddnusEwTD0Ub2FsIYK8FPgO2+zKz5bfwM5wHaR
nnpcoew1nUbhWEuYxVP1lBspFt7zgxgaZupKtxSDwN1Um8eYQHU4I9eRtNVnst1ugOwO1VEZc4uS
WUqQXHYpUD3oKbaBgFBK/Co58t2erlUIzl3+fc01CFi0pxsKjR6TBX+lzdrpZG/ySWokRLdF3lnU
HIcr8P0J0t7eMGRme/WbSZQBvf99+LKWjN3XZRZjc6DsAiBdSlut7qBCDqITFTZQwibLv8m4jyyP
vOJvwIWyQP1yfg2SZFyoSM70xv3iyxYtTWA1DEXoWPJbZzNO1BQuPQo8RbhZyWshAK31dLgVJu2j
UuZt8TRtlpHaAMGQAnrGDU5SCK9YGI1TOUjaKHGF8Hpo/QJ/J54+HZ4UXmwYqkudaArAzNNlledn
0veb9B8cEaudATOVZ2yJmozruVewLL6/0eg+JdUKagC5yVuj+MgS6apxUejO4kFZZexuJHQbcMWv
SrIfnpE18DSamQd6ODtGrD1sxxcTW7Jaei5lQKQIzAfutnxZffAyctJot7DZh9lzAkH3clu48eQc
LfI40ZeFOJtjAyvtfuGYl0AJHpoZke/fQnAWDS+GgUUB2KT+hm37DKxBvMpp24JlZkjXtxbvH7ld
MXu/IqfCPSRd7vYwhQAq3PXJFycNYzsoujfof/qnlZa+sCrprfLTCYC9B+0LQDqcS8hqLo0o3NSO
SVZb4IkajalAk2evgfJ3n4bs7Mk1gIVCnYegcT9lZ4ouc/PmM/Rnhcj3yMRUUJ4YDfNajBGMnvVI
s+IeSXqZ5/yVqe8ZyOCYujiLuxjfqHEZMCK59sph50nqblelJUgHYzvKsGNQ5ThqI5XCjKUos4l3
UxqrrZZty/3GpjXi3hXCJY7jyxpbG7qQk0L7p9HJA9rpcp4DZcRtXZpMdVVLvaPjxsvzYRbXOKcA
qNIpECT5+k61tdqyNgozmwdJCa990s4NIPraeZY1zEirYWx13SIzWtWPH/jWuuT1spqsYvV7E81a
TjM3aTKtiDx7TIHPiIvddBb1GGUxRgmvopFOTHNBnLP/1wNTMYlfjZ0jjoVFaZvj/hFjfAwQWNOF
wX/PR/39QM02x5fiIj/IE1iY6d+zH5OWmYxPZ9AbkRPAlGMfS3Yxtoxs29H0H3D5PvxTfAY1kZJh
9ZRabnjAnuKLVZJGz9gtFKsQunS9LPkHQ68BYcmGxTpKlbCsWAxZ6R5L3LDjPsD0AdUJqm4r18DD
Xx1xux6SpuxP53CgkX+ERxOCd0YjTwVGZ0vbHfD7WrB8tNv6HIcFZHk8wPdG/BAehwlmSBZAwTra
SsfXR3xxFAsBaQI0VtPgbCjFPUEy6lqM/7M+bV6MckPWBc1yk5J1nPnY1ewmo8GtGQQh5ijJMSpB
X7fsB8PFx5IdtQFC00Y5f8vTuj2jPzjnJ97RV/eUXDQ4GrizlYY4T1RwYyG8KYcvOy0McA2eWgub
0YN7I7GDLlOv3XXtpDoYs/sUllli7GQW7MEOk8/yJYPyvFF6/nnUfioxvQRqIotVjai306Zrg2ie
oOnscbPi1MI3dALBbEiarTWimajOQdZXiJZv3knS1qWfa5VxA6kTLkJ3eTj2l2s+/77ejDg3akZO
oFTZmNFO2kWCYPKNCUY6bvPKCydUSUpnS9NMEHvwIJ1HW4lcJnodQuh1bxFbydFC2BW/Xiq8YbBC
QeOqrqE2+RuwcRZRuDw6K6fKJubpsnuZScbh84x//rY81Ca5YPg8JMGn3uxCF5yQtwGXH9My1sXh
/E/Bik4NBdqr7cNnM+w/PBYBpmoTMTq8KiLDheFbEGixMWhnaBxhet1HSQmU/0bYVFXxpyZoHUVR
loh1GcNWvT5cJMurEbB+n2ZY79B1RG8JSj/vpCKJu2ZoSbH4hCRTicELgx9gKNiDZ4gpaftteaQu
0k8pe6GC7eMIIUWeTcChZPG576D3rzx0D/Vn+U1TU8OsZ3JWz5RmEmPePAJQDZSt6kosafi4Dqd+
G3A6uQph2o4YcKzL6rmzjzXdITl4xS53zuEN2rZskfD9TsTcYX/mP419kLWoxjslCDNjen6nOp28
2Xv2zSWh7oXJiXXrRD7KAkhEEXsm29buSsAtPPs0WMddm6xdTOHQg4nKQYUIJ8rJg2x8ydT/Wy9h
SkklmYTXRyaAmQ0gzGFtZxYH91lgTeCJiqI1BhACQWKmvDLZv9YYb/n1SYrHnSxDA+QyYrg74iCv
5VcVAY1zUokuLrDtkoGQ/7x1RirIdMRPEKYUyFhb9xh7BgqlZ8hZ6opTDBK20sHuj/Sd6iiMhcUK
Jwl3BsJ5N0N6uR01D6mgSo6TA1T0PhHQu9fycNs5mGIAxBz5FXSOuIfPhnyarv0MnIEhHw++jD28
q8wdffjsKJF+PGM+q4lIRfMv0vOWkAKDLXb+zt86RWkUQTfQX4gumTIdeYm7EbXiAxFIZRkpsUjx
04auj5wyB0LBnlFIWn9j70HdI4WXlQmi3goVNtityGSH5lWdjiPkC4ctTMUhS+u0jDYplsihARZv
VDyDIubvrYK47cac9SJNIxgHgEiCeaYnCT5VEdBbeY1fj7p8ueSqW5RP7U1rF2piy/9liPpEwJDP
chIPz92ise6h6dl1LinbJYWhSBE1JwkZvwH79aSnYH8jetDQ4zO9sYa4lWLGiZMUArephfye3m3B
1XGi1eA0OIxrcSdQuIQgwYFqTHXF3R2fzkqnlN246sgwMv34XyfDlZ3YK7/dclmFET+9TDxOhKRF
AW924PylvvKmpKcboz/Hhr6yijbB6b3MdrxjttpY3NQMjg00AwcyeUXMR/DMe7R3DOBZ1dMVbbg3
kkHDdxT90iSkkcq64BQ9FF7QlgwbnBB57cfqoOqOCRujd0JDPxdL7t757qGIk32WE/62nZcUvzEr
b+fVd4UevvrDlScQvmZO9zUgMR9oFnJZ1P3gkhIr4u9e4SPZO2iic3V5wXftaRGfT4dzsrZ8cmzr
W5E0Qcx8CT9SbMGLj6xgTRDWrN/WXB/IQkYyCmpu0Z5DgZxvm/A1THS3s65/0ttLA7iQn03CbKe9
Cios9CWjzVeah5DwOr8NMHR7prI5N3hXtp25PdqaggSSGDV+As/uVItYYZuYaPChgM+XkH9lUsmF
E3jzX2O5keFPh3uMYAydITg33o70QbUhhg8lLSlpvxTO1HW5W2zMz8+TEkKV4K5QzHh1BXu4hk3M
3txL/rQ52d+wxfNKqG2bG6yn9VXP3JTbJqOPvCCAycmvVuYokXq9llE3Co1QeXzSki8vs3Mxt99j
peOFBfa1nImFaF64wVa36KAMU/5aZvfiwtvWxvdngPqXO/P7dXqTFX0PgEQ9fN/66IWJXV1EltAP
+RIWcuItfNmozjm9pZSph05eGTbTYnW0RSXhXPerPh5LbbiMiSBxiAOVzM3iJPP4s3fpxPLHfx8g
jCu41xF6PBQW99e4MEeXLyNkobDPVnT3/o85jxdDmooDhgcuG9scCX4GfsnTfNs+bzcQE0x0XzSR
rdeP5l6PaXvBrNpyndcOoTCb1KsTz4QkFUwEJk7NU62qmkgPWDUA39O4ROQoowzUd1UBHeutlqHB
uDccDRfMfaWQ9E8mkvrUOW29C4sfyguT6RryvE4+QbV7vHx04fMDcwLfwUI7jotG6dllZJxcXIB0
/412NmCNV7Kd5oa/lGfHwsQo7CcAFhsJuiIi4NzusULzIPAyeWDvuNfri9kmZuIe9sLaPS82lTUo
FUun7BM9r4+PyPLDy0k7mUgtWubQ+sqyT+RK9/jQa9k/woaziHJcxnh0ApP/lvbX7PsSrOzwlmZf
w5vGHMm4sbSQEdcGgbAQpQ2Wfx05kbBTTCiMu5dau+RxpP/zlZjfd1JIo4WAqu96O19rl/s1b1hg
+aAQXbEFndPU9kAsR1Z7KpOXGDDYBRV9r6ro/lyLI1rNcj58+svQdAegn8242H3dCQlBJ4Lhlvo+
TUnZehpuTPFMv5CRev0aw1YhhEsJLV6gNkyAsJ3qLN5uXAYVvtrNENh7a50DUDw5xw4GC53WuhV/
q/Qh99h4cL7ag3OzpWa2YmPz5/Z5DXUaAO4PVqfuijM751lWoqNKHLvC+vl2CGc/z96+cGB53Y/0
J07IxlpFkBEbsMulf/jrrqUZtArSPCQ5RxR3qr4kA8vCA/cJ9NhRKvYC3eXDh7eUtk6b0UXkJ91V
tUEnyDKWVYj4oig9JGQJvE3alD2URMuAyCPw4ci6r/eAq/XNM3PTxCjFe3SqwfQvV6BsJ/cWWP63
0ZZqSbRbXKa/6wSmyqgU6fW4yb2MI0624pzbMrDnscf/xC6UgJAlI9q34ovXtY1Htp67b9bEBdpS
AcYWkd8lydm6jqgHQQKZdJ6r8H6oei4I4SB8zpoCbSogoSXVulwLaIpQNFBUWyluCXxF3ROT0/NX
da7aXPkwTENlrSdMexPApvxY5CfS6ZhosDieSH/8c4brQMbKBynPIqdj6m9k8Y6x68j24K1K9JJ0
dxNSpBjxJwtU6rrhw6v6hiOnHqvd37xCzPklLNnVUUNHHrv5dfGWgXHgd5HAXJA8biRLY/nOGJOr
Oxd8CYkvblBZsAqXelsrbl4oiMx/1dGW9KJFTGKgJ9TM95EuXfzDUoYGmK7EFCBnhFzklIHTk+1s
mqcqCAcLdw50ZPJyAU9RoyOlJRpkPqjli/5jduZfnXDY6D2LFq4vmhbkYwFHEjrus2VVq4hZMlea
4ix5YezTtw01YT1B6S7INZrkyfHd3j/z/kp4xQ46Bbz6lNI1jLqPsi5pzxJa+ufA8JCt+JG12dfF
+XWBAdbdDD1tl/MjA3ljDioo9oXNC4VTA+22svqPXMJQIqo6VveH0DrsFstkxahFwLKyX/8PSXZV
MlccUqutUarJZELwZcH8R99Y6WY/yE+J97XLcp6aicoIdEYF6BBZjnB0rTY2mccklEEkjBrjgF5T
YWWgnWq7ffjhWVYrB9BaHd7QMAXoEUg7V7glZufnJkZeSOpbJ8ejuvdnTDpexLXORZjessoINZQF
00Y6xkC40hxQv5blq8wgzAH+1+MOcbLg4ymc1LMApCiXiSMALwWaPGrc7gqK7bc9kcM79uIByZKh
tnmiF0WJ4FsFWGeAW1JO0XLnrD+7Z9b6GYLU5zDxw9GjgcyAE9Ps49kEek5buBafqOlmrH4LoCFY
vZu3z7H0lmmbAaMkpfDEcuZT87w76wXJcGJp3mGv8prTEYz9NR3CzKpBSfcD5zSv0R49I9fBuXs/
mEHZWUAlpwVlfShIeVeb19OHb6Ug638Wvd4zOl2nu8vqQqaGAGDQpExTLxCXq5CTx7Tx0dhYIb39
IKQ3DvBGxzfLJAVESAmyYakewSW1F3Au0QsAD5K8R+ikVNELtOenGDQOUTPafAPgZDyMh1QiZyM1
M2nlA1LNHpebDZk7QdIxxz3KzQHRCJkybwVa7duz1pIGdmmCw+lIb2ZwNQkxWecf7U24iWCSPfsZ
cRha8IwPC7MjoFq0D98CTyPGhJCgAgu1SCvX2nBCfTfgwVsR5vYTwwYuGirzLcMLOJ6mSZbQvAGW
4xdwt7dWTSO37PbPvXZCBC46TJKl6MgI2tpm7RNx9M5jKdTDsMzKn8kB+xtYAO2OPGGoiea6rqHk
RjlTKi0AIx9IL0F8GUI5yd43zLzmDjL10r/9FvlxamsB/+6I4vzL1N9LHujHHALTwoEZV0cxo6cm
naUGNZjP4WduBpX5dzSWOsTMa5usArWk/SLUAszX4ppAwynGuIGT5DRVGAFCFY/9VzVXIryWqnM3
iC6IqgeqkHxrXaaRr3fUKNUcP+geUHz1kXRz8K33S/gM2vlwjiY34cIx29JwOsgZ4hK+icfL8b9T
S9wxd8xoDaWBvf4d/jZGuU0cyGFjtnFS3VdIMrfyvmkfm+1jrqUqrKuh2gglHINaos5QVH0SDSTi
tfL1kDH+KA2mZNJ1PDM/uWT+IfvUyPan0g/3iKHXFBaZs1+tbKmUf1ySfXyY4R8Gxtu0eB585Ng1
qrM/WgG/5IEGH4ozkEGEWSMjGqPtTGUkJElZ+gSUa7yWOQjoL8jlPt/zr5Rw/BckyDp86tLImoPn
3bwtEchiMGmRw+GhhMmeDN0gxxPcjjggJgqGFPx94AeKVEFWDiko4TCWRyVGaxCLyESF5s3xVurp
uYEupbCuHt27OYMa9+wcG/gfpUD5QGQGPBTxKaeCUWB42CF94cMroG585chEr/YNgeEulQt1O2i+
Iz5C2Unmn/s39YeZBNsOwAISQyvlyNqd4RMTVgt8Do46b5uorqCbFLGYA4EzCX7TeSO1yBnxyH07
edct7pCsKA0BKTJDFkWeS5IAQT4ENLJ3BsmMOwgPShLm4Wxh7goM1xKQAh5G7tmGE7KeY2MdIK5a
jgL9PE6fpuGDdDOIsiC5M8pyusDQGDVb1CWWZiFM2sl9enIJd2bj0KKsriJxN/1X7055gfXOFKUp
wUkkKkI/Lwp2yhq6/7VJPBkfr/EJtZWvRcfiSdr/M4JKYTF52nwIExf4INBifLxHF0UnNJPdG/VB
ehYbT+eFyxHpXkyvkzm+st5vJhGJVSG/NypBUqqPDNVfptAR3/iVRkDtPpXqIrYfAquy+qTFeu8g
D7FXU4C8RHUZmHMzSh8TaAKNt2wY4qLY8P4K6lXciPEcPKeBtgwiM9BA1teptezVgvdDRGiyB7Pv
gdiO5N9newu6vj0Q1gFJBKV4A57OXoZ4k3YkXTmbkS6zEvqiizFAOhzheHI22P+PviCj5igCJyhQ
JHtGZBVUoqnfSohT4czJUEpc7XgcB6+Imt42sudHoIL0SE1hKsXimtl8q2XDhAPHfk22AWSY6VMd
6f9GtOdmn2c+Dd+UXe1FH6pMugbzz4Z9LvALr+sHYBLrjMH2jkvnUn4kyjZHQHNwd2ez2iVMZy1w
4Wlooqxa0dR/gSOSVo6sPFS0wBxJYenl/ujl5Yf1IgMuQrxS6lgVGYDK3UtKO7jI8ebt+FPxv7GQ
ThLFwI2ZrZlxhKRfOMgp545Rt2wsQQtu+OMSB9MJhD98sB6Dx1ZG08yj6/DNIENGsmm0D9O/ZCdy
bTzs36k/mRWgrl2N/ZxDCrTV81Tv5AuPH51UAcaiD+TAOAb/y3M55HKa8o+3hJZ3Hb2rrsBidKVS
2CNP+cUOm0M+tW9wJuE5azh0YDYdJU1JNHWGZR14zC8vXimSKG85COnzUUFpCi2dWb4zhnjJsFBS
C4iIuSpHiYEyOJMdt9lADBt91Vw/F/ta8b4KVSyzRIeDJMryeg4SmHBpBI04609rbpX0BzE4nPr5
aCTFOL/lpZ+QG6sIa/88maOnJx+8pgkCNkrKneQ2XIJD9FJSDViDfnzOpujPM0IPoZRuwIaiDI1a
zH1PpFt/q7B8vCVQ2Pi7CmctnAkH+FOZQmP/0fkqJFSpS4qFaF1LhKZbZhtVpT+NdVVUSNfaoo7c
g55svUjo1t9ImxccKVAWqZbznC5YnCMBsGortchb6WRL1Vbz6RuGVsWKn5ek+xNX85kJo9G8g8vj
XABccQqC7q5EvbGu9gepqK44rtDRYKCn1s6ESnVNs/QtcBbjBoZDXj3zVgWhBTYtyvRY+IwO/rKz
nIzvCneehfRYxOJARLzBo3gfoj3fEgRP1+OOYDVCI1eIhXhMCaeeNiQoy4Du5+QzJxVM3LaoHCLe
P30VBtsKWI9r0m0hMGS2DRT5O3CH2BN+JFmdho1D5ITJdQKTEYGclY9P6FeFg2fpb1W90qD+7pA/
syvmvvKiRR6LnLOOs2fmH3Mp9HGGFmsPT2RRL3gDnl6HJPY2lvpWt+DLJ0b+6spTPHnGms+I6ZQ1
Rz97RgWCZRd62RqVoXTMXke5G732lbaNHHQN2GAHRmNmtQGOn5mj6ErCofa28RJJXhHQDqVE9FX9
ajrvULyv+YLlM3xQH2zHjZMYfkiLo6pDnWawQKopq1sD74X+uH1BbFl56ITc+EDSHHcG/Qf5WjUF
ZM0TMZSEmCaWyQd8I90pYGBuG0i1NSUaEwwx/yMlvo77S7SZJ0Df4ppbox+IlUoDjRsahkt3O16N
lZO79gX7Q3CS72mLHDiiTdZUqcgQxKJDi5Ja7WNWWQi9j95ev8QX3ma7O4dRPdilO/nZRcAIx/yo
Ce/e2//t4ouOD8aC8v1rEMonIUTdL6XYDFBV+DdKMk5h+PI0Bk3ftECHcmSyWzFMhg2Jjd76A4PL
aAKbfrtVSinNRWo4XwPKr/7fuGDsp1s3mm5BUbdD8rVTTifZn/2Gnq2HgWGBvjuPAZ/F35DP/Qzv
Y1AbMyU5GF7inraSfAyffw0fYeuaXE8iBmIIXn7uE6Fhv392OGlhwDROPKIyO8wVFMgCuFyfecq1
Ks63WoyIJhMcjYNzVyIIhk1yK4NoEQlEEkGH2OyoUZWvRs3JPPwlJL3LNrInHRhYtU43Mw2hkcJW
2/9Or81Sm0SAFYR9Tuk/2NQwLQ+13NlyLK2FyTLZ3Wn3ImRxJPJ76BOtSrD5ZT1PUGP17ZqPgWf+
QBJfkJZGJnreh8XHHdi4UvfbAASW0XxjAJksUmGkmdkfBwStijYKYitF0g/AI2DE4CFy/yFCoUM3
ogdegPXek3JlUXJboVgWF+O+dzChA4vEKhjWuVzSx6RjcIl5EUaDWFsa/wCCB8X08/vE/OQWAfcE
GTWJbqVwBJJQIZh0FNXJtC59njosMJaXLMAm4l0E++icHAA0Dvp6f245Y3nqPrSGC3woJgquICd4
bTdN+jbFF23U1k1MNAXG9XMo6dvIw4A/TVdVpQdk8VSqfNCW+8l7MQv/SDJUIpUW/wKVLdNZGY1p
5ApDOkQHFEn3jVV8XR9ck0rm9+dj9LtqZqp+yo9wcGSxVKSGLjH9VNvxuD3akIFeDRxCu2R7Wnx1
MEfYN6KuIvU+4eOqkecBdaVHco214IB5TIBFbhvYpGOEoUenIKHuK2w5+yEErjlzvzdaHHY0zK6m
obtRwIINVxsAHgwivojm+6rkjfiLREEEZT1Ux53slNWevr75IYwO9hzytBaIAvGSqrNQfGoXnXmK
9wovje1G7I1TNhVLKH1m2//AUdzgYleo83LWybTZgsaOIGb9FuoRYKznRhAQygBinQeJrkyEtEnz
pvNHOovryKTeISd31o0b3qHXHMiTeysm2m6v4HV3GXYeiprLMAse+POtPdX2CktG9OVFRIIN88Qx
EI/Iii6F7vPMku4Vjxi2LeFJNk9JcFJkvE0P4zVq5kPIQrQAQopyY3bq/v7cl1A++2N37VK+oqRo
rGi2n+/ip/TX16WjwAwB6+eJ31oKEsb2YsSTk0BhkmyP8a0i8UlGGJBJ8G5AV3j4JKTRX1T4sMBF
pe1dhJcHgRM6F5Xtk4BMPDKgQ1+g30a7ZWLPgDv4w0XZ9ddfGfAiWOPut3kQ3/F2XU39x2XExuYC
JpY8ZnSD1lrpYVJbtOz7RRSP5sRUCnuOVr25hZ3XXnVM+j4BjvDKnt0M2nhAca82TgTSupvcxPYa
y0DiacKCx7bjPUnWRIlpGg0Q710OKA6uVOA1ODgEkM1v6KQ2+t3JRaW2dpClDiRkEzgb6JFJD8RT
kRQ53ViPYvkBS4AoSoBMt62Z3bcbDP2mqzqpSLcPbeaQ6tKonfjDTzoDXRaszXT8ATLgamXfeu2n
5xbHgmzqtnM2Z8k3l4B1G7iTQOFU3DsrcDNyrGqLz4K0BaI/JhLxEo9GPl9/SVS2ctl6R9B9fSNB
UXWeUSunT8ylAxCzfumW6SkQ8SAnoeSdOOj56QFCgUw2x2SpYOi/YTvo5HkzGtY5hjipEGDaDrlp
YMMKSWp1EaucmFTecD72qOmzPl9xZGQhP3oBYfJG6XZjypfNuMAYwct/O5JZc+RjN5L2+kiu+kAo
iu95g0Lpf+WwiX7UqAh/lwBJKMJwL8NLE7Inu5ZrEA1djK4yr7Rv4Pkw8xmqWqxG+wMbVit/9he7
nqtDgwFYhv4I0T3aYplx0lR2eoCsqnXol22NrG6+DB3kq7iLZufxUIlXSMyVNt+H5DnZeSKCvy3T
0Mu1cAsn+I3VxyCCIEVcRbyRYe9Ftw8MTDduO8f96HbbMjgcgaYPztT8aW7KUtcJKGAbVAj3JRwO
b4ENW7n4QIhT9jbm9Fq3MwNeYn5+RCOQjzkO3kuwDdne6tqpwcMhVpCvJ10bS7B/r0cPy9xI7/6x
N5EEkl0H9012BJKo3k9nIeHePrQTevSb9vcd5rvsInxU3PLKyZ7X3Xo2FA8ZZWdfoshYDENET4MV
NPdZIvl1BmGyQALj6T3JYQ+STseKVRvieRYQrtVvzK1OyoWoJT2drgnM4nZzgEc8JMx/RCyOuUKj
WqI/eq3XMO1kXFMpvsK1vDArN8pRrGp+ENsWxDrDBVgU1VPozPwT3qvJO/wOkMiJjr9dBvi4+rKk
o6M5kzdSmYPEq9f840gjJw8TXxBExhsMHfE02lsGQRtTLA2mY7AFqTBvrgLFSfQzwl8Cgn/E8kLH
swwv79/xkVNVQ3IgXVpiWe2rHBOSYd0e22toioiTTXXywe12dakSjUc5hNNWg6rZnFggiHqW0icn
WZL0lU6X2M25UckZ0MzmfiwZZxqN4uU398+vsV5+bqCs8TMFFTyBFLVZIw6nwmMJSozVpvZB0M+W
aX2BrM/GpKQ3GS4bPs7NUdgwJqVl0gePxuFk/hw7m3L3R4GKm3WgSUXsc1OIKMtJmXsRu3iizZst
xKUlW3QNJTlWBgHWZGJh6shrIxe3IBeS/FA44C2eis2wNrh+Wj13ilxaTFk2zxc7TmU3S5cowqQF
k/Tqkz11t2aljb9X+81SMW7DgJMWKPJimxaNCUklINz0siL0bUN9DEtseO8ry0DbiNApIPUvSLWX
BqlIWD1xdZhhV45SR4qdLhAVcJssiZjoeSXXtNEMGLwFsLCeXEW8EQocZ7fXlkfwhZJ3s5+Jq8Zz
46c4QdcDCIFgcfjpNlMQP8wiNSC7Y5VDw/7iGoqoDvy3XpbL0BwICMDjauIWolUgUsgcyh/ODOBv
OEjub/OfswbLNXQQoYQUUGRXrIQ0EaUw3pApW6bf4jJT/0smzvAZ+xt1qL7+kVS4IYCd0QNfWsiF
z8jKmtf5EK/WeLmyd+lyoEGEOI2rYFD1gKHJ8b8CG0r1BC3D6ZExHjetA5TFUpt/CVZeMLZR2zg/
ElEIChP8CtWOxYF0Tg2zSxkkYw9hDYppW26M/ucBhZqx5fqjY0Vf3L0lZCO+ptHUhCj0i9ssqwkZ
f3Ixf9VzaaZ6dfPLQ3F8ueZ3EyeoaFMIVm0akNJno78N+EmosGcEfdnC/1u3ICCInLl4BqgP5yTd
XbKwVgSnoJm3BDvv9BdoSXSd1c0tU2jpXObGfYkZtlsUnQNPVFGTXDv2Qs2Jb/HyZa883hc8MBJD
QcxES82dk2ammi4i7uHg3E7njkOVOfVU+XpzG026e0OFETO0xePfyayeU+gJzIc5/uSxQog+Zoeq
ESZQQUx+5hkTkxeyr/QvGGgdMPhKhzstSFXkaskPM3RQPqK4cPCmJaO3jG8Sp7/NwQW/u9hjPeTc
XMVqYVntyqvXMXFF0p1UiejlyjYoFWfgmHOAkMETkwc33iP6lt6tcnYn6FHy1YVRQvJpZy0aKnHv
OxvYNUKgDmb2Mey+ppAoo28lh3JD+8oiakuODmfD7D92QFc668yyY3YjN8cLfkgp5PRrw3CbVS7p
W0BdMNbV4c4w9I4oQ2U3rS4nAOYyn993OgHt7/d7hEeWBylOc4RLCaLAafN0unQCmVlbZL7ba1mN
9Mr9zh/V48tZ/I4TpVGWR1rNmt9C490CNrOM1kQBnv+cLOkuZFQVK3EJW6XkMEv8s51adYZpOnuM
i/ENA07UPI3XEi054fyGjwhRLbF4IyN7V7oX1Hlm1sjB3rYts+/FIboUx1UiVgXG/9cwd5BW0RAC
tP6G3JkLnzzTLg218ypL8BshB0BuggtbSCG0HnxN7fz9Jf8Jc8JNPQ5O1kJPB5U+K25rTtwjWqum
Kg86Ll0YlQTHLEsRo9fRnpZgQJG82TcOSS7xih1dvWqriX89LrJ9omGtq/Rj2+Ynxdw0v9GFUTH0
XCgdPQLce8/Rgv4uCqJDnCrHQyXkuX39e62aDB97v4VzV883n2YN/Ti6s6DPsDx7yCYrYMAEppPX
Uh5juWcPDlaNM8sD9qtwGYsfLiwrniP+5Q+9r0mpHez62Phyzfag13uWSkgeNGFH/k/WBRZTKbBA
Q/pO8soXP+ScIkTgiIPRoECY4+QvmqzV91IO5xKuII0FlB9pnVqtygMslWVgBuX2aoRRhWBZwjBa
qLn3ODFrBJqvP8o5pLKGY2KnPZD1DUE07RaLyeXqH18LFK8T2E5hpPz+eB5f2X4dXJFGY4CF4eEd
t5mxdHToppuhdS45At7msoPHCY+XgGJbVEWmD8LHRReKoz7RE6dxeJq17/ZdeSTlWx79W+K1sWic
YCYZqzPAYk+gGTlI+Jl5rKq6sThg7n+FIaeuO9SshZPZlsZ16pg0kkxaQ/xWm94YxmQFBA1Suw0u
OR0FxNVyPZmJWO5IVU7jnYmKczvkMCwA5C/QPauHeopj0ZOokOXt/cTKaHzzNj8L0qfpjA7ltMFi
rB2sjAqpC+KeqkmyzVpmE7/+OUJUTlj+0v7pHGlxbl3BGkc5Wn2I8fj1hWMixDNAQL/6QXVBrlm4
nDwlwVuigw/xhVFpTTwFCFakHA2Se4LvTKgF/n3WWj/+yIthkeANzPBC1o/a4gecy2JweTC6fQr0
ETW03NiFLHU4vczyfYzanNMm8k9ymdTHNymx0GIxLRVDDdgRBOM8RgUjfp0j+uG7em8sngb0+S4S
QEahPOf+CMO10tQT3+8gH23ALQ2uHiUZHy2+wwboo2gJHer3U6VKwROx5XTiNCGuJTdti1XrCy0P
mr2MhTxyx81etLKJBRqCU/RgNIFTKVegLpELss9MC3G4Xfeha94sTBpYfq57G3475enW43kDInvy
9TlH1kOwtdznHmPH4oC6W/TCMP+rSe5t2g/qMY4ZeLiBN0s3qmt4x6DWVni3W0c2Wjgjrx5S/jzx
MGwMysCobOuAtb57GAfHebC5DVh67miLX6glbb860qo09wpaJLd6GJM6ZCpTSuXzaJyOv7H/ti/S
+/bYiya6GNTmp8Z9+k5AsDlUM1XqYPYh9mu8wvmgcKu7xd46KpniivzlfEqrUzUmc6fz+MWx/vmo
nP+VyzYU+dah9smcAwCPZw/0DcPWb0vjXVNzLLN742YQtRlIsZXClqKP0cME/67QiXlZt9l9G/Ib
VXX3kmT9q6ZvwH/vXEPLDlpLsVraoi2eEN1fd1JrnEhoezElO9OcBsOCxHjbCPP3ZuOeW4Ub7QVl
3CBgNCj66IklfOzlI/7LcQkNJE+LobzL9DET4gqfwcQR43XU08KvrqOiC7SX8gcznvCDxCpsHI9y
WQrtGSsIfnpfHfk52VahLwzpIn2Q9W7e7KlIeN3tbaCWSy4OUPkCHy79UVOg0uZXlgLn4JB2EvJi
Ap266MrK9QQW/cFVx5CpvoVSsRIfu2zs7eIPI4oqyyzWchPYB3W0yvUa0d/uM1wVRPIdondDoHEz
WEtyecwFJfGDuqQdYz/OaPb+IDCrcXJDQIDCme5Qf501yDUjhyIfSmJEeKkWAX2GHBSIXqHqtIaO
hmh4UhIF8W8GcbAFZdwEMlT0lq1yLN30NuApcDMgYSysY4AXuK9h3zzX6FSziA38d8Yim4HtK/Wb
5xwf5zrR5eB/eHll+AWRSr+1t4Cu5TaEnkaGckh3M6jbLKRm4TpX9/cPXeF6wpRzdF1GP/mWaEjw
qeDMuvksGslhy7RQOZLU8kBOhA98lcENVxvwYMlcO/oVx/kgTZX4k0w/ImPvH5OT9yerAAwfFeM7
eBAMQi8zeyhpSNFUrpp7PwBKFymY4ZC/XLorvnQF5DHWY/g+g9wy3QuVNypK82+aeMWBZdD7cxff
o4S+V+YWKOo3MnC5T8ov/p2dhnkwV8e8/9NiEeuJGgKEId5oBkVQI9fNFQf13cLHRZft2vhnp7mT
2Mn99jmQ5y2OCJqCkXuED956DlVwW0yqAEmBdnE2Ty7fVaJCGm7h3jhy61D4IRv+SdGio+CxeISC
2cwgeC2Er3+/Clj1dTRsYZHP0g8EvDE0rGQQKLfB8FcvqFCCiwij2sdIJBrCBBQmgPg+Zknaiktz
2pePLoHwVAZ9RMWki9ZchbOOJLP+uFKneIwvZv/+2zmul3pSuSgYjjGsMnp4lpjJz1KI0cDRM6Gk
uhK5uV9PgH9zi85y7oW4KzZQbxlev3ZhehSK9PoxC/vS0+qBTiPRXwH5gb4DHXJwVNyv4n7VC7xX
b9oPrgevUM3yxqtpIfzxay5Nz3kIJDJ/7M9qrirL8oXhWOH/zpKMKdzvPPjOc8gJJ64iINpqYIAA
iwUljwnNT4dgJRnNYHVoKp7zv5xpkW608CfDhtw5/8j+8FSV8Oq85D1i/GID0OuP5rbP78ZmgPKJ
xJmRpxjL4+hOmfIVaG9q4A3KUnVn+zdpRr4KqDE+eQO/kaZ6JD37MHvhzNFei9i9swTmsaSvHvQn
m4RvjkM62pG9bjekC9XMUs8vLHtDGTI2Ab55l2CPz9sd313yQ+wTD1+XggWgBnPv0E7qilFcgVXx
5PGpaERYJs54RzpKUGwN8nnjLWU6pqRqgLYseasie9O/xHY5ExFFKVlNXSM3Mog3tU52Zui88mpF
lETftVUmS6UIk4t5oYxkPAZUEIfHonmTSaCudDQnXpyz2NVab8nrqG7IpBd5+uLUfLO75DRbcdfO
jCyO0D4B877Z9rR5Q/I/XVMoPCqGqlNN0fueSslW3DSluycJkHltDPr9Bkbuzj+Pcowt5fvPXB/r
Gb15wJExZ8ayEy/vJfag1v0kxaQfY2pUe0oUr0TsZaipVLvFEhE5G2C3tfbyoreH5RewdJnNpvI4
u1eL6UksFa0PVvqGTJsGnADZJ3AXPFkRIaLBFZZbmqzNAx7QsJpKbNedyijZCPCs2K1y1t2Esb53
Jj4+s3cQ2tExuPANEI2aTt+5M8kpvjoEGJ8KiaFQ6edIDllDsl9LaqHoFCwjryf1yX8c57Da29nL
fAj9RnTp231RaJp2f7xOXRUHEkJ5Q0xzDNJlkE0Ue+lBNLDlRpr7fyLTRiCiYuoI0pvec4G/ZIBg
S+8LyuULWGffEp2iNMpmI96VHqBWjp3mKA6KnF4EGyF1SpI3iomZFuxWpRnTk9rVjuVYAFOtYLU0
RBFPZq7Ny9Mdhlo+nYS+qzHubrGFFZRY19ScleR9uoUuNhuqq0zLcQ/KAref/gZ1xCu2OBhjXeto
G1b+MMKo+sjPgwA5mx+22D7F9fkToHkoPBefX4G3QXJ8ozeaC/u9sLHlFVYZv+h3wrAJ+frH8C+W
XsT7opG91PjB5AYFA1/FtG/piVgxrBxsXwTlmfleljaKbe+JDt1/DhzYoJL4AKpHq5N0UiDWQ14P
iS3LtXmyt/yYcTchFhjmE+4ygcBmkhd8fOzoKV9WkeVgr/UO6iSs8D19KXGKSgqdU497CFgIlPA/
4WjSFtNE2m/V2RGzuUKYxes8KCE3LdCzf+K6uhmlQD/r4lhpgLgCVby1Huw40j0fgkReaJyU18Rw
AOyApUC0IiFKFdgNd97mOY0VJXRRYAiKQ0zc+Ppk5ZBEvLnvggLYxeeT7/GasJTdr00I/Oly4a17
WTRAhMb4wtW1ZZT0LVn6/wkupirRDaqDIVQiXzyenPPF/VvJWn5baepeKAZSOdjP7FZHWSn7Koji
8C4O4Rkjz3TaJhEKAhWY4HUd7O1Q/BHGbqOwS2K7TQ3woa7ytAzRanDn9m3Lz27QEwRlcSATyJep
zx2uVvUil3RWXMHvNxeToNf5jEyeomRnWznF3ajVatnetOnaf+SsgcuBFdRJxttbT3SjisLKH5+e
w0VYYOnHvm6wJRyG4JnoRIByGWR1eHyBUfUvrTJ/WUnBZrxUJ5iLFqDDGxomvv87tzIrWut7Fv1F
1KGUf1wucnUIxqaiQKbrXaySvZ4pJU38fFWD+s6NBJrYb/i0VIH+kdf4p9MPWqmUlpqmc+7FSq0j
6eSLDRGr/d7AxDKC5H9o+rvhTkWbKiiMuV5aUK2wfKgKsaIy6yCP6UWaT8x5igagmaHK/xRNweeI
4bfn8gHEcxif3Rn4NnlOLv8O0lcCUZiuvqGDsFQCw+30Qx/Ykauj5rAf9RdmDNoOXyTZp54Skf6V
QI3Gn3ryFgXEx1msa3v9iU6C6Ve1SfNJ5Dmaq3/f2zgJze/GPLVj3Cbg3qXqIaP5OGbgCqv9qvVb
NccSb6w3KTyfEZRGgyuRsKXVSUGpdmbz2nRUxMGPaVyrb0OyDEDlHQScARuIQSMPP76sAr6fpIzg
WZKr7XibusI1KjO+BibwbpMXvh+1wfAqvTMDDE+NvK8hYRQwLD/e7zDPfWx+OrDky9c2dZi2bah6
rDh6NLlJDecbd0d2aH+LvVMB8CdyiWty96cqjuUpSEsSe2/xnQTncWMFU/yPiHyqXjCnxB8ZJ9F6
DnallDZEWjC56Fj3ZkQg7PBzOPERdBzDXJNVQh4CpRZvrcU6TYZYOsCJE+NidmEFib7xWRf+8xdj
QlbR7Qr4xYe0to1XX98gOjFtQzX4d4uQEoY13VMZyafsL24at4tjcsQjr680XjlBPiA4FwjMC8w3
Qx7L/9U5+n6sH5TqBeL6yWtlajZOyF5vjtyIFScZgh2oj3TmVXWzPmSheSS3yIh/vVtJw0s3TH6g
2DsVKW6CrKhHqKOxbkQYsbtT4h4AW53+ZuULsX25N3Izn/ZUGE+s7JiWhmn5hK0hXRc02HF+6SSW
rIwPvQoGDbYvrggl0exRgNM5fDKDwFIXMT/EDDf2wpnrrHeWCw106wNsZEOgx/vgAUAlhf1b2sx9
P1mzU40RucLrmumO2OH0lfrxOWYELFle/gqx+PwkGRPTKuZDcr1xbtPth2x4xH9j40A96dqejOhL
Mdf0CO3zHUKO62GKXaCJjOLCn0EbzSQGNHyiXPUJOrAOgf6LSaPmHyVfTspTZXpw48RjzJ9sK8ji
DLwNHOZ7wMsu+gZpiYjOuHyvOEUE6CcXl48mBp7lI3AnorTrZ20FwBoYps8K2PhWMDYEUP+CKVSq
CQ+p4TrE7tskRb+5B3+Ata1pyd+eUbe4Tqg9ciQ1pkNbQYaDHfB7GNPz47g7YhW20+0b+5dhKRM7
ISG/PGtX7kOPUfWFB/WSNVenmpdJhaXonxyR71Y5WN+vSgD10HdQc9dn/CgLXoJyrBin7T63BvGp
rutFn9WqHDkLRQJGlo5nXxp4enJ7agErhnrSa36UZs+JLY/j5tZg/ouGrzoa2MFyZKKC7nC1VkJJ
RS3sNYyKhv2Wntrr4CUfQgk/zchs1KlpycxbFnSHCQuCHSmGFhNIrIJKsAQqvBcSGsPfnS7ivyrQ
DIIqMJQB11GcavjV+IEdqH87UAVVH3w9rf1BCzV1az9p9Bxqeaqo1MjZ9jZ2WhqcQMqraTPqFCXp
c2hmhv03XwV3ofL3LSQ13B208fcFrh0ZlkLhSj8yO/lueR+MSu9pYuAe3El1qPQy17R1Xe1Blev5
Z4X6ixS+wzeyW2lSevb9OMwG359FB0pL7rHy4rGf9RyMLYt4YBiPSLOuYkkPhUsaT7SaqMc7gUHM
WLJxicInJV7t4L5er3/8fzd9IcjVcSruYwd7TIOiAIfU5ctqiMjP8vhG/UBNT8wSlP+RzhTiMtxU
UU67Rgsfn7cvMQ+gmj9+jroLKXqkbD8Qe3PiE0LlmDozY8A3NsijgxR3ak6nkqyO77mYYBK40fVr
1BU9/KyQQT245Qvi7JNcNxd1u6ioueOFJmjsnG7hhcai5Yxo1u8TF8WRqPrwJVTz4YR56a5a5Ktu
44f/UDPbupNpCfLqPKLmyeRQxdMvifqajqwEUbW9csTwXzprfzMQJS/0IquBijFJFFApH3d4itDh
Iqn2dwhDcMlxDbSNLBDvgO6Syx0803H1InBU8oqnpxMkNSWQJR8RD8qHCu5B6Q7pnLB4spZvGAlY
EdOFC8ItEfSVLtR/dqKeHC7GNqg08wFwuP8qbfp+YQxh7EW7Z2lbCshbDjqa4QmT356Fk8H1qGEv
3QAJTJCtdiAW6oC0T67gzhCdNdNcA5IMoRWL9vsCUco1o0VXLmB5HQOzW5Pld1d5SVkoqmlwmm/x
7ZYXKNT79qhkoZ28nFfNi8CCFiKieW5zPyEb4wlfkYJM2m0OckHDqlRckr/ga8jlf81OoIEjr1Rv
GpCHsn5YlWMT1MijsXiT0S8Ki/iL9woMziKLayHg2vsTf+jEQuffv4KWMeXScT8vTrBxn/ROPPgZ
x40tNzyvUR7V7mvlpYpCpeIRC4uu4I0KaW6+7rtI2UpgkXrkLXZ4ZSn6+lEFwplLVYXFY50o+iX4
YQYT6UNkhzQbc1edIUAMcm5VXhZLIhW5GyRYq8K54kXCdF2NJ8jQDkEVaonsA5Wysfd9STsjxVr7
3QZSyOQmqQKeo3mjqBq5++V3kC5OA/lSFJ+uU0zmWyykg3jsWRbDTpRCrhajlHeLjDHeIlvg7gFF
qyveUCkiP2SOgXMF78STBIIVr4XiUFn6t1frTZDJv6bArNMuMIroes0Mmo6crdXbWqstN0SgURWh
c3Eo+F8kS+b4g8/Sh60sfWJeQ2yH4Qz3MtUxBtgALeGIG+pwjizEDT0zLtpXIHtWRAAI8hvnMepo
kN4Hv1G8NfqrvRpCZRxXgzcQFJqJOZhR6+LcMDRmL8JyWzdEhborpXrtv11vwMTJ8T/a8K+d3JHu
kLBFqx5S6EhCvgbe1GVsYmkQDiyWwqNAH5y2I+/hSoJgixxAQ1k1OZ/V6PDAx2Db07O2mJcZZpub
85lSz2B1LT+KkWYY2SaXi++Y+R1NHI2mvUIn01A+p/qgIzEIkUNwasaKi2D6wsXBl2MjartHLi6p
kkHQ/RYnpq+qs3xFXen/E7DBidXfGGJ5IFMkBr3YzAGmz4Ya1fm4v4JAeX0jIQszJU/cuTPkkfxX
a7FpFBPmjqKwyS7YXLSekwHRmOUTCZ3+FhYBzb3E8Id2fFA3JAUsC8spnf6M9vkL+k+BLB/+tTUA
f0RqVzQi9erpzC0HF4Rz37+43WkTdgPdzTwrSpdaH8044YS79tttvWK005pkom2lnbajl8tGMlNg
mVThbQz3GSB+EaHyodriutVEppT08lwvv5CgT/yVFIfihNO/kK98MU8udL9OspGK4N6iczt9ruKm
CVnayGWbbYJLdwjDT19wtuCpOmYbwbEE/qggbk5S+Q19r7Qcmx60+DxkgrzZqhoyZHHOgsKMDsBS
39P1k/ZCKAWVISg+9Ap1cyoEGsUApUp5KLH+fcHS47a/mS1g1GPItIdSL0xk7pE3P3ZnhIZ4DtxK
/cQj51uaoEg5GS51LA1PnOFjjXYupumhRYTbZo3sDcQOli3c+KNrGW6iJB/592bSg75WCSvaBtxI
b91ZJ0pZeuaBTuN/Z4A82AoYS54th73sOQp4zYQqbbwEovdxtuknAIo+ThGZlw/LGiA4u5pciUAO
UWKNWCTTZcHenttE8DCxZzHhp7R+iRZ8kokrxJYg2us/bTiKP1VKQNVqu4Hp0uemss9Bq8GQOmKR
cG1FRU76uz701W2hVwIAjXZ/eqegMUy7iykYHv1LGU0yC7nQEbsuMIVrhDB9JulwedlMhCH1zTRn
8W9riRHGF9Xl+ahql9lm1LOFkJ6GbhaPRVvS5wVHvF1wd1AX1hcU8hLlTcKZZX2XfQXiAl5t8s9Q
ym0OI6hdNanDr3S7m0xVoYk+UGbxk1A2Y18WfUL9iJz13t8SAAILmtTAS2AtO/Moa00Fi5ZdzVU/
RIAnNkkOywcEG1m5mWtzdTTH1OulusgL7Kndp1TR4TBS33XFHBnjRVUHAzDramiiwzAIsdTxO8yY
4wqr/AZMw9QPA+DOmlApuTOjQM41WtPS042oj5icVUaWKD9szCJvsVas4Nn5QgEwJMZiBmAlFB1X
SbQeuVlSVnsbp34ZdW0ZKojDxuILzXzCXPaKIG+vTYgoSL9yOrRTBbdl20EXZyog2TC+xQM3X399
Tn2C+Kys9v97NkNdS9LTAVAe7DmBIcrQH3x0OguuJXNl54JYzjv8LZaH/b6pBNL0lqmjvzlDRIAz
0jaazC//MmPjoua+m3dFL1omlGWbKrzoZ4nhvtw8BG/QGanxPrVNVADeNaovJxkNF+YuYn22aEXQ
u7/VILQm58rX6DUGlDah0MuuXFfRjplgnFcYm7bAxql+o04u69cLCZ05mtV4qYZmfhOXQeuRG7fO
nOBpZ8J1aOu+/VHJ1J7cgpsXheD2agJHT+ttf1+BhnvvFhv6/xdIHQYmotw3JFxs5dFAmS/Wy9em
XtVT7tV8MVT29s/hrztmjqaVqPtUGqXJaxViqRsF8eEC6X/sBKRLV+Wf7OzouK1YrahaocdHyKi1
wFvb2zNU0uYIOpNaaajHeK4HIExLKzAJxheE9NNnpOvdpiJxl4Dm5A4domcfvK3wx+vyAbd1u10z
2u+DNKBV2sKcsIsXaVEvRdlNK4R1ndWbSPcxOFXqJTslJGbWJbSNbII0Kr6OO+sxHChktcqLN9k0
HMybsKrhDTfjYy+tstVKCUC9BCGqMRtW1x3cmWePbtEpiULhhBtEK0njnLRGDehSkEvQfyBnUbyK
K7bpipQGsVY6rSULrqKBW7wflejN9cFb8j7wZjLMjFE7YV2E+pviOmbGTfcxcg3tEvrupbSBvOil
210ddG4LK1Wsk4imxYYPb4zBOXHBZDft12wjq9AX16Wzx7X1RpoH6MXtFsKTNJOACQP7Pss97L+R
8+rRge0CgdNHY15drXRiTpHWa54Zqa/XqyVFU+tQVbjPtzakPn3fteveI9RpKcBwa1YDoVNzBR44
6XOyf6zkpEwFLXJFiqaSc85lbxRRvWSdFsLGyttnLZ5PgbgqvaaQ7vqbEXcyFTW64mWurDmW71rM
B/PPI7QyHZw1sjpvgPWkaIvsJE+Ow++47MO1L5nbkFi3V7cuPTa9wHhGIjR5UkBRH8vkmAzm+E3g
XsIHbCLtLQTvVQMs90nZ0mEiBs4fRGelTuSqF1rBpY5vrlG8TcwL5YLpW70ud3VAE43cnwRetSHZ
SrGp+5/fmIC3Gy5h6CeRZs4heMw/Zpy3v21dqjDOImgXGiZ7GeJmE+nBPAl0ky8MD1XWV8G0WMHY
e18IE8908CwjG8JaYgEkr02jlFhesuMCea9DaUyU/RlzK+KeLgmLKFUnmkI3KMSrHff+HOrU0grk
6SzeHhn0sNoIcru6phFUW1CGlPYkwHRFNBA+L9Q5ou4CgPB3Ka+paBTeunQU7tdglmclqm4Gvftk
2ZQpiRFQkjJrWucwBGfnMCD6KyV3N7vhJZQCWsSbXKrhJern5ngjJh1UcLQvxUb6TsbBGEOXMcZ2
367dZMk7jKd9wMVDyAEtCZGsYBnPRGSADvz9WR0DpYBTiD6l9fJL1/aN9GETthLExhZjQFYb47My
jDpMH87hhOjabcuAgV/bHy3lumaT5g/OV/yRTvtxohUoEGdpXFlrokD+Hz2iL6CghJ6EVfpq4EDw
b2raF2dNh3vGWJKupS7ZqXKUnHd9+dGvrYOhx2Q8OTg61XUu+Wy727P34wvSaFmBsSOtMpBeGu3J
qCbhxi0D+o3FxGrr0nkuYxDcc3rPUlLo2yQzKlGrdOEQbR+ewY2TzlMjipedwUgk+EArdY9StEPm
qckD21t8ehMDjXx+SE9va60M3a4Uf8baOEKf7qib09RMIZC1UxFcss+aiIvHi4/zbmZGxookB8u/
iI4Y2QQ7CEHatrX967IeHVDG5bBuPWT9MzoX4dJEy2Z4dikurvnoSkgiJIEWYV4dwioIg1izJl+l
wMwAZH1cVYzhZH8mhbCf6yJfQjCObknhigmnSTs+KFJwJNT/YN5pW3As4hae19sqH/WaUukAD378
KTL6JjlebwfAx8cy6Sc+7gHO0OFPK5iqGFM2eY2DQLtFJ4ujA3E2adeFqSRfgtbyUv4atO1t0Pwm
Gp8g8R0Xdq6rUCus+hdq3peVo84LgvUvr3MCN598BrCp77ojhUim1G6qaZJ+cy2Sj0KYG0COiyT0
hDdRlS1m13lCeZhNmgKKJ2mEU+BftalYuSpwatbMabyMAbIU5KGJjE3REaTR6Ld7FC0k7dkSBgOx
WOC7jfANCJWehL84fGdWBA5nrxu9jYA4yP6MrT2eDRB6TGzQQjYfrljjGBqkf8Nse5FQWdLgdsn9
S9x1dO/ZgptKh2nf6rgYVOafkR3Dqg/BsuuYwneFXB72P2AFikW23zW1SzM294wQOJI5dHn3Fh+M
nsI8pv3HsxgRoTTGlUUUf0mNJPJ3RK/XHhlB5RepOCwlDMK9FUqBgKXeOx62y4OOvyS5uYjUPqYb
J3cBtpnprxEKupZOlQbb3UkNH+5t1bo+TI+mUI0idiIrxgP95/CYHF0Scz509/9EichKKPFJDH5u
1pY3cA1A5+sii6P6kdY7+7kr1zBp6vGnBRUd+5WPT78H/z34UNhlpWFt9+lXaTil9V80Inf3qlSE
oeTgNdE03uiCg2AFAb5sqMoJ4ylWiVB361Pnpl8tXFKTyhwEklphzHa0TtXfZh0LwH3+LPzwXF6q
OO9dulN0JTOXv/YQJpfCjQhX4fmhuoQhHubd40bx1XruVkm2UY1m4T08YbKuQXpyaBx9siCVoMNR
duAm13AdGM6tN0IDat6elYBJbdq+appr3OyFce/oLo1gMe1GUJQ3ftnJU5Q1uqHOuhJSrpY0h2m+
2TjJS/WVpur7TIvIsm1jh81YNWq7bC+ADV7IsBZsvB+jdjN7rDRHODVgN2P5mx8ZoCSJ0o8MyjJ5
axgEEWKqS3hPMpQfXM9hn2x0X4BgU6SuHSOKUm/2+nscjOaZKwqH3SR73/x3gQNZ3hNgrOUT0VBA
fc51Jzyjn8jYZ85bUSR2rnSiR2Osufhuvln2B0GqCxCikIc/czBHzK+rNQlKkLhmS2o2jYmP1l/6
vH6DTmfZn5v6cpQi7hi7DZ+pIgE3XZOPA2wJtFs81ZtHH5E+83QM2KheG1kpIJDVM384eLZg60fn
6T56j/8wUJ0tg6AvWv5gn52Zw2jYiZLd7heieWX/PuCOO2dy8iHUO2jjt6XELk5g4nOHtKj13HM2
8Gnd4HEVWtWxIatfHB1RoDBuQzMFukLltSdNGzHXuiyQmZjEuOOIf70uHWtRqy8H+fPehpVzvqlc
RaJRW6zsK7Vy1hJoe0Nh00aD00s0bYshYSV+YE+KGgiZXn7OAVggs3MMfGDb++LRn434xI2Mug9g
Q8dS2YWBaPw+L87S/B/92JxiToUSrgVvqxmubNF/myEN/KwaQjT8tfcN18mF2zo1PgXy/1A8a15M
nNCLUUXEmdb8ZIWpfI7iizQc1bsgQXRsGjW1NH/CPvGz9H4kBFcyZM2C87rLyBZrd3he51XoEuH9
yL/6z9LLaXzeVmPGR57Ecwz8w+HhocKzphLlSp4YfPuzTj/4HScQGmBJeZqmR5tYwSF9R+Qa/r56
t7rLkQXVAQHp6mzHwwxrOgrBcZU4taYfKRphP+dVb94evpFKcU3THI+xyeVVZ49CrIzqW7r4JnHN
jhymxxYM01g2T//sRwbxZ5xgKiTQxjIJ6uYskQBeNY+SiDlLtOWMmdzsJz1xmXdSljGWSyCnGsCV
jZar5XcNvrTi0Hfh+B9ktNos6ysVMX9TQpzsvjr805PpxScgw+20UMZBlAXp9v0CebTBB5KUQWvK
c5uA24FOumKQ9C1FobDDUsvmx5JgLal1VPSMU26j8RBaHWCrO/4N7xugywYHlUwMBZCYD67nKQFf
rfV9kN+uKGePqSZKunWHCd346EzkwBls+hQ1t3RpdnJxJIuQIUkGKuxMno0VNWMxKkeX3Ef6uNp5
3LE5MNcwXxd6STm/G5gDfaqm8T00QWJ38EMPeupjVsEzwFrajjxXOxEFM/4As6cxNR/yd1HMsAk9
LCXJmipEit5MD3VTPDYn+LeCscq5vRJIdtW22/zIWChtihmoA79cXSHID/YxClaDBTKRMn5+ukPj
5ZdVD/TTg24aZwz3BqQ1opY3EOtOv8THZ6mNVzLnvKhYvPx+3BU7mZAUMx2jkfrAX7EwAKhv4PuN
zj+P+lZi1w7VcD14wjViuSVOIq3l509hdx+Y0AJJ4sm5tX0agwPK4elNVmC0vwpD+oTdGTkuxD9n
3GV3bQPuJlF9gMWfeZZmJI9oC3Puu5QIexsRRTMOJoMr+KYZaFNeYINTYKpicefciy/IZZ15ync7
NYacz1Bb9Lx5qgxCnHHv0TEhq/ip7hj/wzz89rTWP+sTt62qedEfyHSbv/lfXpkaLsGpAkCmWcjX
1+WuzMCsXsicocUDKbifHB/w2WUKryQ32RRnzj1TfOgk1TbgKoPWE2qvxUatT+8Z2VeZOh5RzDGL
UJOvh1PFbAZeozaWouh30VTBTqMvTXyyeZ5MBXchprsElH5ucf7ZnEgkgOu1HcSQwKVwTfJrm+CY
QFW+rCqJjJMBXxI49hhIOrTyMewv3knovax5TLMC8qfj1UcggFZ0MEx4OaOKHFx4UJGosymVBtI3
Oh2xQL2JXyw0P1VYXVeW7d/mvkwAgyAZdfYYIKA6u4WgdqBR5GjLk192zXjocAKyGl6e3+14oCZ1
JSzVXcfk2Wy2envyryi91pCi8DNQJvBBP9AsQLoL5/ULdtVnqbiC1hRjQRXZfqtpVuAoaF0OTPj6
9fEN1grfkyejmRiqZKTH103CTg3kSOwRJv37oIJm9detwCtxrdNgRYdHShspuIRNhAQLhEvP+bMR
QGHTs/PcNCqbB5M21DTKGUnCQSQsYty3XdY1Z0fbyUu5r5Uf5HyOkpjyQ+xHj/X8EOVxYIWR6sFx
uVhL55Qpf9iCdwBvbyV3WWdmO/NJVv8AQeHl6fzJpBBb+g6yQJhdgj3nY7tIcuY9L2qsDlM6j6T0
h2x+yuNQt/HiKZp/QQbXM4WJW5mgEnJEGIqLl4gD9NYVauW4VrKeez43ifzPOUEF8esfF2Yv/F0F
14lr3/NPUpUROfFuZsPHAWzTfeMfqTI988PxBEAu8FCBVQ8mq2DH7A4J/1j8k4jITi425D+A1jLl
RTSyRgih+TDJm1J7U3K4d6qpC543Urr6ZhTcAEhYz13RM6zK4PfQCMTskj2fJF818oPvvvhI+agy
FWUbZ5t2vzDgG9LcIVYlllGVV+TScOt82pX+ThNzc/juN9m/so23F13GFuLDSti4tSjVZ+weaxqg
epaGL21m/k3L+K2zhZHfdX92YE3MvHCXhB3SwhRZZgO/dIxjyao0/a4Ue7MYWlB+BLWVkCZ7rYGO
GyasZdcwat2tYb9uO+bGslJD3vptPdR7bpkkKxLCc5C4nsyEwtH/PMftwV/VO03HFwFsS0G3/RQf
8HWl3ZPhaosx14Sp3Y0ih2JgNCvcZCjARPq63BPih8US1XDGuYJCrzKeq8vuwRBlUxI+2VrdPhOe
oRtK47aQUw3vW34mAVH1znBpvAfGa3w3g+89RLoUGSFypkdln7PuYfvPFlJP1sS267BJ2Qcp9J7+
CGcFC6ypI7HYpMOS4EAd0bkgHkfoW1ln1tnhfKMlEZbN8/aYo+ebWAd2hHn1W+KMmuJNAzvdWsHd
VZ9Br046OxVasaq7iyRZ6XbHjLDTqZjC7EQ2MGkUlMqXAvBLreN4eITHjaKUM2R1XhzdXfdsSxMe
Pg9yor1Rv3bo4U1qgxc5r24nrShln0pyMyfK+sApUoPaTgyAN7qtJ1LSkvDBI01YngYnURqnG45C
0JMLgIcMaHzkme7Q3U39n1fSqnZnn/AQOAnnxYGZUfcdZY5R3PG7NySsRUezsjTmhoxLkyks9u4w
FOXHJ3DhUJS3RdxKibPI9vfiWir8WVdAO2803QoSw9c/I36/pacs2+coEZWvz6iAJKAu7EQDZpVo
x6qoxGqN2JX39dGOpnlBeV+HRwHRKsBuRoEpsCgRc28o0DIBf81rFXFK1hitzE88dohfh8JXyv9j
2mMfUz13iRhT6hAvkA8vlEaYBYdkxdB9m1qH1+2RreO1JGSbnbfQ1huDDLpsyBL8VDJCrzVGQIKo
V+6jxxTTC/qIZyUuscJhfl1o0sE+SKdsT+fHmI6GHKAOciYypqUnAo7OsIBCEiT6e+KhD8cO/jdb
DvLk0++ezaaULZOx+Lede5OgoMPUOsMY5l7Xi9ptMh91LeCQCHhxuDT73xx2elxgxf5F0bVx6zKm
NC3AMFBfiVvFv/i8C9Cq1+DL0S6pdCq9zLAsmUwVBuTu8di6jxqKncCuPLCoDHiPnRtnx7jnpmEi
O81LoA3P7RuITIGBeo9d0milPIXJGMhC3SQNd8tkri4KWUSSIr01gRXGCMnP4Xht3h2I6+eBgi/B
ZjY7vEXdxmq0sSnOcTo4CgoYcQBaDuk1l86YfsvJzu1eBtMLyuQzUQqaIDEro+JmG0Pa8Qn+HJQo
ngzRqg/J3aDeSBJKpJ3HY6sLOGuJzAwSWrY6Ad6qZA8lfF1cG9zJ21/Vc8Wc0z+e3EGoVHV7caVG
Q02KC3rUrwohdqm1GxqgVQ0+hQc1XQ7p6XlfoQrVsrS84OXvydWHfu8QBfE0SFPhjGYWLk41a6gW
a5+/8FRsy6WzWQZMOg/ImRruELIQOdshTeCTdNxzDQ4HQ/sylTfP0944uBi/a6Ywo81APoPhUzCC
F0FIgA/DVaRf5DbZCvizFNgv/LibPZTYYDeL5WjIW3PBVc14N8nX5WP8BTHTUZr+0eCjrIhMAAlS
os+J96DA2wI8m2PlE4YlN3rSmehJ9qy1HJbMGLcTpBlfwBwF+fAxzOP054LwEYKb3X1muuNTJUG5
PkfGOD6vFb/ENnNvdyaA/VNuSkUKZ1/6kN2fLCbQuwSiV5M1cFeTydsB2Ag/UpKWG1aANAfnyxU4
wpBKdHxTlIOfQxyNWC4E4rw5cpq9ycEBo852TStuagljRQcJvTkt7v1u5O3OMDCWgo0Z0V4FMcoU
AT/uNjXmWI2EBjNgDMcp/Nq81DKqZKq+ZfY54iMWRo0llZ6VNJ5BiUoprTkh7p+gX4FU/jgVDRHm
JgagBZCYQImWLksrNdV+dqhA7kOIBWLRdYsMfw5rV95PNHl+isYj2FJUwtTzkMk4mW6FbQ1gpsom
Udw6RuCvYMvblOjfowmHERY5RMZeDskwihkHAcQh0llgprzaV07VViYuOGFVUq/W3sAM0BOuco8l
3rHqXYTLM7NIhI7AuEfboFibHwqsJ4gA7Hr7zFIkFl9QOvPjJBdKG8Xz0d+RorMYcHweQJAXMDXp
KIiScROF1p1uxtFx0jz+L7172Rl8PZ07rt2swTGS8KKdtNESUMAlBquT6MRpBSUxOz9iI71UcBqL
GoimwCk3jXduxIi48cM6MBDKXG0pKQj5TvM2Qrc07diFviNY/P00gOIGXVpbGUQG1ZFs6MCB289n
WlXKZSh2qKAJWTW/5hIrdHGUoc8Rz2u1uzYl7p/P22mryplcBKoxu8+ryDwA/86qOIcrdJ96RbPU
jqL3rkOnmeuFXUThmht7kUM7+L1+F00q5SjD74sYS6w0r1wiVmABLSfnWWk1Zc7pZv/VgRY5QbMi
WeGwfCTl2+NuS687w3BANANh5vnSYgeVYgpTjJruencYKSEYHkKyQsXvti7qvKEu7svjkzL6O355
5EETaEWJ0lBaS+WzJ8TbYI6RLgZXRZgtMwJ4LmgEqcj9qSc8eTvv0iqJsHzi+Wc5W9V/1f/M1ke1
vVRM9KLfyn8Wc6fDriC+mvtGrqx/9zXFaCGG2/6RyB1MNnHnxxD7Qqf/bVtPSUkZEhB1vcT2zGIR
PA0+XmFRsjUFpVQz/yH0O7I8Jog3NxWjN1ldXo7UxGozHXgCwf2aBHRsyBJd+OKbuJ6M6+bnpBYW
KQE61lZ1EmSIGbHhEDYH97NcdO3SEop91336yDXTwuULh6bpY88bpAqYCr1aq5xNfNisFmeNdCD5
CBClYzMCwYkDPcd81PYZ4D4exg210SzA4UhNkqt7gsBY+C6TLYESmWVIrL8plfTUmSRjEW+Fb/o6
e43ZCX5c+tKx5Pu3OLIe4YdDate4iPItAV6ix7jq0wLBcMCPmYPIJykvZ+wGasDWyPHnI2BrL2m8
+sZPOt4/SVvsUX1Rrus0McLHbThjRfvweUqetOC+zQ2LGEaaBHHOpbCxauZ9KMxnPlI0Zmxm/poE
3EmoLfSaxa+dlLRtCUPxV3fhlTHr8+pnHJPI7E52QCn9TsC6r5qiCsBYCB3uZWr6cuNA69yIsnwS
Zu13LGFqAO+QWOVKBOgqKSfqA2PPhTJf2oGZ7r34q0SGEJDvpP0qh7K8FsNeLr76YBvQaLg5MvrY
uqClRlg7SVXO2SIKUTXiibj5bJW3kM8MpEIKLbf5d1KqvOB6cQPDhMEXEjtQhOiQf1gTWTyoWn+r
ZpiY2noRJqH83ZnNTSV5AlTrVSNwrW5mJ9sR7tL4ZXEMlenYAUc1h9W16n3SYivLcSdJXuX8ZO59
3UGauU8AndktYVLV3xHLy4Aw6+X4qCU15p/6X9+oaubQr9WbKdfcA3d7WLiPtMf5S2D5dae84x3J
nadQCWYj1gq8/mvph5uWbxB3usyZ6Hl4lOWD1u0t/M5wryQzFZ24bgZusR8NZlE8RN+vrhXc8XNA
Fy1hNF8j7oBo4E3AUt9Lq1mY+O0hFJoYJIPuup+M2tbDFB+nNJqBvkWFMFIafw2Nj6tsP5EG6dKs
BUtDZI5JlykZyJfGWl3dOeukrKR16rqHUFGH5BKn+/b2Urv+wlhdfrsb0gvrXgUEuFVbijPx63Yt
DxsoUQEIqwK2PEclDavQh0+DckbM30hLhmFiSPk0xgIiYXgCU1+GP5+jHMC99oJZXbfNnnYR8wP9
2UX2PlNfv/tZgHoIHeQ3Gn+iq5wHe6BILWHwPsUJS9TUeko4jszjCeRp/HHTpCBDiwHoy1dgBTRv
2i6Yyasb01GEN/qN72i0CXfmCEv6ivEdlgD8SSg8RMfKmX0kg6/+04WMJ+F2CMdT1+KgvIEDBZN+
AqXrpjDW9KyvoHUDr3PuxHCW7uhlC7B1stfvMF5N1qCMc4LdzEW3E6Dn7OEVTpM6G9X+id894PJ0
AaFL0GNTvKO8kVZB+N3JSoefF6C/y3Mlx69IM2LXefrWaqprXbxmWMTgTTQDhcVFQ2isHkZB2bDJ
ckRw6EcqSgLVJfs2mK/4JKsVFGAhhmmMlH/1gYTkDI4hVBdHlV7cjNSlPN1VGKJpLLPKtnN8fPys
FXQlerZWVk7WZFDUqAJUD6QRcg5C3lDDujJQ8XNUw7t6lwjqnb1+2ZkyyofmxniwvlCvxQSEZp7k
v6zsxERN6GIJsczWwsy4CUej2i/ClwkKELoZyAt380Fu6nRZCOi8Qp5uni0fn+Jl0pNxKBd+xxEb
vrWgi1lEOgnciQRhgbG99vb/R8P6iXQS0ipc6EnVix0Dq6oR4w6YY1allWorgWVYn8vrgiwuDm/V
RQu4vz3CgM4gXHC2EbsC3FKWJlS2TgPxCE89J4nT3RcpmL4Ghpz2rxGHQV+ftQno1Nw11WaKVN3F
1d5v8McOe7VH8/Y/e4QIUv0NEFzDUY0SpARRfEIjYO8ClVTOzkzsQ3c8j+BbQ1IRu1IbydNGihIr
LklZy69r0X/bFtZ2qQ4CHIxpO1c7EKXyarkat6sPs46TMXAIJunsgYMx5uLrLeosCJ8QZT+xA1Lx
t8Jxh1svjqMI1kd8g5YTJGA5HlBJEO8zFbn1WdRgB1kRsST1g+oLFrREFsEzFnfPOSt3/2XJa9rx
9msJQ3Cs6l7DHNcoP8Dve0Jt6rwiguNstK+SYAUU8reTw9XolIj1i9Aj3WlssEo+Dp5RPuxLBtH2
CvXfXtL21vMFuGIgfttbQQbZPEfHsCcf+BSs2wUCI7OfDN/BOIWnNAUY+kjqIBC3HXGU8yUl9dIN
lFYC5D3296OOvXPpypY3the0K+hPVkRnfd67RjwPdsTbNSuAIPykPHxQu6+8c48LTsDCMHoyyt1I
i7P6ZtCmt6SE+3Od/iMhkqsAbAhIUeO5f/JGrysCf21cRKZFhZZv0TX9MTFis0MfBUDdOVRn+6bb
HaRNMn6c4GG7wdj/oTI4mm0ECfx+Vk8kg/7/2QnRAJvITvDF8ND1dAFPZopDDWKiQNGay3ugZDjZ
0fk7XSz++KiH6+NreUXj64WedroII6YmWSXV+PxQKP1icN+CDHoDCNJt1VtyrcNRX9uHZ4Qwr0ax
L5MbTxJvYLYPPxTMCB9Rl8aHKUvSgXiW7z9+e1cwvoPxKCW5baT/9ZqxcYHEG17lyb7ltSpCm3Kd
j8IoUcN+TRzzHXspKiwWe1h2Il/4Er9yrzitqR7GRkuND+/evqSdSjQGvN9C5XC5huafhC0Jqfuh
arjo9yYfm+i4vQUv4AYHRqoKs7dYT1zOPY11DbSf2MiIghRlu6SgpuAlG8oYhDqlJhpInIR/9DpJ
h/qux0isvJtWvQOC+zdLiwFtsSJeOgMrJzUBlIIWHI0ybayXBPwdIdXdGo37fbVUZiimDxgZKeWd
6C1GsJkNL1TWK81K7YnG4ZNeHTyhVqT84BA1/ji3qBtopeJY0VTPp8ov5NVGbILGPhzd9jJIO8lB
S8xeW6mFneDWwA/Cye79uPNrSBOTJ1xfC0fzJbIRIu70K0wRpjom1FcDKa3O8P8tYErXoZGdY+9k
zF3/HN9ZP7xeMPzDJFySPdRmY76pCWb8ixCzg8F/hLckkP62S7gczivjdhhFa/Mw48Q2qa9vr2/e
ilITh+M0WokWaamD5Qhb87aZSYEC6khUVYhX6dYDh6l4RKLe4wLyxO5FVLvrOCH/p9X5yDfp2h21
kNGefbn9hvGrJnjtJO3lO5rxZBnBT3EfSdXtRct7iysOyg9hOs4Xe9chBEWXAzMuL4eBpjZs75C5
JUK4ikgsLowY+gq99hwqHUjfNe5KNarRLLBO/o6HoOVoRGbBUK2gu86WYkDTGoEgRgKxFc6O43mC
1RRk4zE6/hUYFOr7GsfKxxvM4k3C16AmyxziJ7PQyMiPvhPd7xlBLNFBKtut3HuFtxhMv0Zc2Hc0
WtJu4/6nw/KlrQRte90d9aZicSeZ41cyP/TMYUjV0WK2IdwgrYuVRmxohPjVrM0CchYG5FXlLQd6
w1vFzuE3ZlAV7cAObJ1m9rb+TIuy21KB0Aym12aPJdhmUrh4l15WBf97Yd9I/BTw6rRr31lBsFGf
fgfQqp8FzZQUWUMHEecrL0cV7+FIR8a3FGoaw6JkxCAVsmcQ9uyWLJCn5bAJ+di2B9ak/iVOGQTl
wP5hp5JzsMqIhGOzg//qBM71JrQlPkUsl0eCKo5UVFMEMRo2ze7vcVRFcCg3Fgku11Vh9LyTZ1Oa
D0+gXJpyIRoUzKjRszKQnfdo+pMHUhP6bsKo3tJXslZ5DP3Zo9MSEIGfNsCAAjt7jEY4AWIpc1uc
huVHm+Ks0U13K94K+Cuq/UrU5Nhf4XX+U7eVS4n0wj+FtNIDig5i0Uc9duPugIuwkDfn8Ua7/8/4
ZJuRVTnu1kJo2n4w8zYJb/5KqFiAZhiDELy+PUgEPe7S3umIGzbJAM69qYWmHiMp4nayVetHNVRa
IJkxNstYPoirPuqhHPaiLeKL3wI6edJuU3hkqondkigUFlSoVRWL4NOutLoF4FPQmB6LUoiO9tlj
exysDb02ddrc4F03OU2oA6ATswaEoJ0oWCtgUud6PzJpj39Y2zK8bdHgr/Gpw24PDi1WIxm2rGMO
mlpa6irb73r3YP1Z2cUpAUIczIIqpxHj4b5egeFTJf2MZwXGlTUpfbtP2psBNMY8mxsX0WjWKGO/
g61H4+qPsGwEH4fpE9wCZJ1g7siDd4cVYukwnQZe9/JOPlpATm/GOP0IN6WkFIvlI8rp3q60Dhxj
ITkwVq3fwUc8hbAln0beKeE3wPwMSwF/Sq3spuhyVWLnvf7oS2bAKZ8yWAUeOSfWtB+gseMAmXYS
d0Z0EPAFJI/VJrkaF84T4vM/x8f73dzRG2yDCr2a7Fd9jggZJJ9cmF9LgvexV0mNzMKsYSM41EY6
qHmZDSMn473Au2dqIzKNCmZwbXBryLrLA1s+J2zD5ALZ13CfB+33nGXHnkh1k3+lWgFPK1SmOS86
/VFN2uw9zv/vLhOAik7J33SoSmOI4QFMm59m5kNMDuojJB96Z3ajiu0Z6ZNpeTMFkaHIhHeL40WL
Lx63BbMTaNXcAA6Z3ESSN2/m/PB9p0QEK+61VotaxoxUB1lIwMd2vKqnl8PDxD7uufay0pBE2os/
KbkkAa39nKlk+qFyc6Pqii0ROMlCN3FKg30WBKfG0nUgo3YShkryWr4E0eVc79cTu1u0N/sTuAXd
p5vYZQu93eJS+jXHhrFs0RmQsyY0lKbyP4U7ySghnG+7yfj/9FKchqbmSGmXIr3M208bSyEibr6+
bXytBtjPFvSItBsjFEkkmXYTqCpLEI67n2nXEvSBRZRLyPWgJvxelgfGGt9Sd5/i8OMSwrYr51sL
4IAxeiEMSHUKLrraHzLqC7EH0KMKozHb/7mYgnjajIuSNoQCt5Ilht8+9HroQrE83JcDwEJBAnfy
UdfulL7HlTuRns/4cLYC324kSCQ3G5pB9Y2tuoNYzaEbOCPpOIA1XO3lnzyWeP9UFwgIlNzQNLiw
kntCjKVq2plF30aL1bKyUlZban0IkYzEBboqu4oVWR4oEkHEfNqWP0mypIHnQ1+9RZkYGoUQ7qfC
eKhYcqCbwhi1NMDBoMFgfvKHk7YZkG8II8mnGnWUvswj0/+rqj7xvqYOUfki7CPJYHfC2ZVv4UUu
fW2lJnshHAYqQZ0MXuVSy30g7qIkpIrCHWRa0Yg2F1sKpFXF3vmVdtleHqhzJCPp7NMol/WTP/WU
Cx2vY0JgiLixPXJVbGuyTdj2IvVGsW7HNB9HHTpY9FG1xDKNeQuqgKO9KptF9AZlUmJx+juFKi3a
10xdz1mAhxGcMaauI1gE2sejZCInzyqrucT9L8Nknj4FDKc4xglr2TmpWk7fktcljGEsugxCA9Bw
HAsYdU7NMeTL1dwB0Z41RuHgIqTCtabdrdEbU0R/9DiZs6err0Z/yW+Avq+PklfYebajFsKWhTNU
lClEsWP0o5I6XSjNxtVM23O1JiQ66Ov6C2ReUNAEO8dYWvcIekZoPWy0duMj8dj/Q8RSGRimZUFU
x65Sontfpv2aiyx4upfhDf+D+rdiK7T5RcFjWyeD6PNCNsI15Di8lNi+0sBjn5A1ymunguphkM2P
YVu7In3PXGCsDtAo+giAJugP6xjq2FVweuIsz628xEPG+TM/FdbtxtAAtLzC3iZRKj8h4/B3dE72
bXaZILnnqIa2zWBKb1vCz++hW4LE0eHsITEVMpeEKtlMjR8tLPGrKO2wDX06dUS5OPZQa20Hdz3J
WcNMqM6TJbJS0FvdsmIqaebeeEtMFHliqoLI229fUAqTYvyYBcAqQMeb0jsDpRSACiNvt6a/w4bW
lLsbaJMuVnvVyUxC5Nkt3Xo0KVzFXLh8el/VAqW2TcZJU4tMpdwAVZTI0lanBnvQlkSgI6EPHlDM
9e7sz2jnbOq73Ox6QdHl3eoE1gZMpvDKEjlFfZxMyc2SCbCMPNRBHRfPkYyif9sMZLhA77yHITtN
d5R1IG+7kBJs4kpiMCu18IWDz7BGAAFlpO0giP3fJ9lz6DY192CMvxja/U8diolwpV07jC53ZDIy
D4wTsVGx7Hl6nwbI/RGmg+YjztKKIEL9tJfuWDt7SzUjtYQAtNKo14lWAlpe7PXe4vazCI0buwRY
5uc9T6s00uS9ti72tv3lzfQOYUbCglKsmKOAB402dEJKgliFaK4TZdD159FsYG2eC2/zj0SlI0w/
HAfEtINO0EwT6y3IywW8ppQI2AG+rOF+jbtjBGngzPvumhZ/gsZZn1bC4uMz/sRxo32vbGgTwVDR
/EPONJ3eBWhzBK5CYIikfRdA/zSOUvSJjS8SMHFFCiZG1tGM4qCNsO+Y0daccYD3rVvJsOEzIJjr
wJGYcKHvlq35zvA5Z0JggexteQGx7J6Ut4231UOCKmIJt/PJZjFKin1SPObCDq0KRi9pgdoCx+VK
G9GCxJ+OQjHIoXTfAM0iOTMA0+QQebPcqUl1YP48ejmI3aUjQ9UodHl4QFJ/5f58ZB9yAXQMN+9E
XpEHUxpGld5HUeEzJrJwMzwjxeXPVJ8RmZTjH+C++7StsSQR6sZ4mHm1j8x9kRIkf8xymwh8mZVz
15oJkqZmiHE139y8Zyzry9QaqCqq0co/szSd+/rXOGFUXl8Kh0loRDdTZNiwdaUVEhQJwvS4mMYZ
1NvfovrL8rj6tq2jz0P18aIQHF5aNKqs7pXzJ0IqY4JqNwA7zVz0tq463P21mUdTeuJLE5oNRntt
Q3uJb1ljYyIxV9NBDc0AixhpyP+iwbYkV20l8yfP6gowuKJ32OVl6O3aRfPgtsFZ8rTvKhf5dAop
uDNDX6qoRoRhsn1L/Nw3PvB8EVmfZDtNQuOr4z7LxFdlLxl1iNjy8RFI9s2Yf1wQpGqRnzs6huxz
8uERpCTrDMGV4uEbJglZm1Ygz1h9k3JDip8Le6VS8FrU6FJNoXbzOAf89bf6GyoLiXpqrEH63J9S
hivSDqtgrmVPZhLfMrymNT7bp7rayuRHbd7V63309sEMtdeHMFmn+tiI4MvDoD9oPKMy9DAgd4hv
jDVqpPsbSh5s8wGLQSRWYJUZ+wUX22NAhbdj8OCgiTJmqBudaODxCAOI2tlJBbZYOBYDM3AI/2tJ
zeKS6a6PADBAcx0p8HPAoqC3MER+x0Cwu7em2iBX0Z/DZucEOAZWivTwOyAdo3QR4oXvs3msjTry
MQDbZszwZF0+svTYjsd/df3sRYkj6YUK1apY8ZlUovowRSPUEtv4PntLpKJsE/BWxVTM4LrpV+MR
2Egknlg/T+ggmWF4VlbfVsJ43DMn3ud5ONr8cDqyWrWtyEJg/S/cKKadPPTZteWXu/9QJ5byzZxQ
IV9sEAvgR88Qq2gtKsCv8JJBYcDLuXRrTjNhtowVeqiiJHK+c/v0SGPYK6y7ugO9mNa0GR89HuqV
Ykdj9a7pwG4UzOwutSiaLHVTZW3XNSELXgcBKC1ZA+p7OAWWjF9QXplIqb/Ty4KTs91/ET+4wUlT
8zLwXBUuSbGNjiTU5ezoBexPcmNwI0fJLb7qNmDvHzBy5JohLCAIWNy92g5fOtuBoGHPSSwzwcQ/
VaZ0WMtc/VeMNlJiRqsh6N9A+/TfzTVmY2e8ry+egv5VIY+Mrt1Q+zyyifLYIx94lr/pHNIBYE+y
ALudfpGD0T9ro1GQb3frDali70AE6olxG9sPF3X8QWFQAKb0mluVy/h5rX38/OEW2q7hXnrbYivG
Hl7n8ExAXaL4ufnakuiaF2m5PC3yI03smL9oPvCkiYmUD6FA0eRXLc5hECZtJuY5SY0+ca9ESLfd
gC9xODw9bIdqpPZ8dZo4OeUCSg/taI7I58fsLKXYLPBFuOm64HrXfblxEyfbEiHlBdGd1/Fz8FqI
f6LAeM+kiX1JWPDGYR5MORjKiim1NPafSllJdgSRSBy2Frih4qLHzq9vmFXtTSkS+oTypyfwIeUj
ZnQpBD9uMVqDycbV8xwr3q+iq0UkMTDtoWIEWyHj8M/UoXg9V/HCDHSbYn9XU6I1e0DJFmIGBDwU
ZXXorQkfNAxcOGFfw/FgMS80+AluJJe/pJbqEyeCKC/10HHJ+dio3YRJvsOFIN8oBBwpVlfh45Fj
qr2UnI3ZE/G+iZJVfcZUyAyZo5qLZKIj6Se0oEPgkQIVZZyhgx9KCDGzdKe8vTiAI1Fv2O0l/eGE
hCu/zd7/8My8gHkgpzTXD1fEferWwUDwAyJulUfWg3650Fz0gpqZyTzj0xRgffdTHSizsrmeMQdi
s+LbJer+0xd4pfAz2ltgfOVU+s03wjF5NoThTYY7ysd/6s58hUEm6Q5SjL+ip2kjEnf+kwpKnWSr
tbbkQKme/nM07vqKmGBhvuwoTcQSzFC2WKF5Uccal6T6024MqW1lIXCqQknO+A/0eQ20yKoBoT8R
0jVPYE+U99Y/nD5A1CrW6cG0ekDOsjLF+rJPUpJDWEPYjDCqeM5k4KL+5MbL8EjuW+CddszyhAsj
giKLnQfkK3aGzF+6sN6Sbr0zYZMBMgBCnK4nrZki/GQoGsFhkLSOmHTEQvmCFDAAQrNvyXMCyPt2
I7zdg3zpyJgsBGAQBPDeUfarSl0ji73MkHLkxrm4WrCkYySKZJsNGquKKEX5WQsFV1vjXW/cxU7h
Yn+ErkxfmLVp0kYOGTZ56JZQYCFtWpQuk7WXWdqrg26lH3chMKBH7p+fqp8C9eR6ATXfjXhd8po+
k/7VcSSW/fNiCiZOHUiuyPn7SDrZPpGSEtE9EeSvBSGng6j5KwFy/4QhEuP+zRnqCDoiQKYoTqjU
2Pelptyfju6y6Op1NRc4jp8ykENDbUhLXDSUS/RhT2uq170sx37dVV0TVttgYqXU5QK2PBeqOUHq
2hkwvSTkRzTyEWaHXUlt0MiWgVlVbzoZwtnjIk1ZriStw8SvBWRjEvy4YpCDqt4n2rEtHHaxkcPN
GHYKgCldd06gLUOJAxH2JEdckPonT9oLBlLBYjs2gykYRt4jftqdEKunrJzUgtEZReYdTulU2T6A
nFiMVGEeGpQR5ZrBxJUqL8XR0pVEQnZ5oXZCw+QDouMwj4Wt/L4LjbMU4qI2zNIG+O+ZiS2YOkCO
yLpWpEibJ33HC5CloLAyATtBFON/41DZ0Y3VFAGd7Yvoa0oz3WyHS+Poe1/Bmlkuo199aqLxw05G
2G8ueioWzyD4Sa7XO3vb9Iqfv5zSD5BzSHMf8O4kKiOwu3J+la6R6OY1h/bsBZ1nAhJRxMHLIw/C
NwDBOMpD+q/s1tEEPjeYboxm1/UgLWcyVZZHxFkND4JWv1VXlFVjFNhfGhgnaxHdzD19xVIgku/y
J7usYpRYgnCSCad4Gsg7k6HVc5V2E3JY8Y1Yn/1jdT6iJRDQeZuNHW9m12JWEEkW8SB9DyIECY7j
Qw8bTD8LXV4XeivNvstM2IaOjpwGRGDDzV9wwJuSBY9saqcHWd4RoThzRQp2T6fBKbZKAQ0mfFhv
SATozOme4H8xKEuYHmZ/WwzMTQCbBS9k/J0hIL/FF55IvlnV0ILdP2WObC8sCvR/Vg2fj+ptsfi8
rcGyTPkV6+DEbT4aYL0+NNAIKO+sBQZB2AZAU4ae0rn0blULJKBQKptuiBcTMZ+jjzBPDJY+oHu/
UHVoDJ/Z4CmaYCk2XU/Sz2LObOgpVoKka98NNLLp2ZFUIGyC7pzPqd1Mx3FyVQUT7EfQOWify61k
LTJY4XT5RRswsPiM43XCxjfQcGUmOf5+prhN8gnGfKjHqo9URtaSHn9mlBZ/ZHLZmrD3uZg1DMQX
z6SZeYItsI/AlcXQuPc2naSNDb6ngat/MwsuPlaKUyejLZrQH1f8Kh5VXYdtTvQvBzfQxDsUHTpb
C/yQf/ZofgZNQ7/Jj3Pvnb19JiIBbgmA7+tCANJDp9q4KsIQo1SQAewpvNXQQZetO4Npi7d7f+LQ
4woQUW/7yNzQdLJoz6VvT5xlFJ28PuDBwOeyZBq2xOcv+DZ2agB87eXO1OsFrKWwtrZyjCW09lPm
uEqGIee7ylmga1PTPA05ptQziPKHNXl2MZkEda3NHJHdrNFo6YQf3X8YPY+O4hLaepzQILDZBYNs
lOmGJXeCXNLBZbUbi8RUGfYyVOn5wL3KDcGrx7Wec1EvpDoskKha8Qy66ZZ6pzCutdWwmWh9ln2j
45Spcy1EgnpoMS0DVbXIZZDhdm30d+ogUxSm7cQ3+yl+WtiPiCySS8ZPIGgn0YNnhcy+BH5ACN0h
Hpyoa5kHF1vnw4NrngdVWzwiZ6Pt5PKGV6Zf5UXrttqROdIYNG8DDX4VMfm6nwYY09dRqdm4HOkP
okiUR0HLvo5b3t9pVB2zoxk5KnRXyGp3cK25BrZoCs+01DtjKXFeMENUEAOwkLxsKl/gozrebkcW
41BrOysoUpnRn1U2e7ukozWRkXbozI3xSoOttAt3vDwVPbTbhzNuBSVxu04MMS+Bo6zx6WonO3hL
0tYi2lW0/6GrFNOkKYRvEzV5+SnzLx6kxTk7ek1wH/kfN42tIEa+EB2BRKFx3UgSUU5iaeQFOFHx
5nSPTxi0mus0Hx74t2lmePCvkVFMOntr6SXRR7tF9T8dLNd4rwQIh14a2h7Z2MqrKt95sZMVS9uN
HKDhkFsuke7l+i4nEYFCqLfBD6xhE3vpUUTs5Sl4hCD0ntypSOwSv8a7NfoVupU0SuXcY8a6zyrK
BM7693CrhKieSYhaPFl1XrS9Q9xIcMSQdhyyPm37tANafIfaYifjsnLWatYa918ByYLjUPOgCo1t
HQZIVdHbGdMFAyvszfclvPkP48sgKAwnmKngEF5tVVo2NczNWneGWgql41QrWQmpBKW9MAQSH8AY
g3X7KfTV+2H21/5/CJjPc6y5uD/VOv9o3WgO9lTEzBVBT0d2CFFw28RmX5BuDjens+J40j4LNFsR
SQ19h7GEovilJkAwj8hVBon7ceIZ6MVNX+Ovar/oTreytA1k2C3UVcTHQC6Xxke2R8tjK722tzF3
PA3Ujov6TiI7bLBL/FHBwGIQ/pCSljPFjPYYdaqcdTlgcnV8zYOBrPsmwlAUxWczA3SUWc4SFBL2
w9biey7k/pT7pRE/zxyItGVifDBla92td5tpgxSSCo6c7xDNHqwSscrgGyJAecjGWU6HE+f42X0Y
cPigYfuvCTnttoU8ZwPJlXlYkPgjtcFlSONHwpZOGtvLi8tPd5rOpJzUDvaE3yQIuaq/Jwjds2Yr
lhNhUPksPcahDDt5zIYKo1k1CokEdC2cqsFCvgy64Pf+0JmwKwXZbmOGVAu4XQVHb9M2PcZ1tc9w
2Ha22wErU5K6lK420tKDl6IZYQEk/mazytHLKZZBHVL9apTtaTAsEySpW0OWLJNeNYfmjGAAmu7J
rtV2yVOqvHIoGkfM4/CvzV3zlZ81QFGxskXTiARiqFEra0ey/tZIgB3eZRPRpqLLs7ZdaOlukagb
kf79prb63fVrqhLSeJ46s2CShUCs884Nlw4NPYs0f9NT44gs9VOmV6TE69eT7Lt6gjNwphzoLN4y
9rM99dEPGyz4jhOjuV8cyhrmq5Hk64SxV7aTA+7YOwVqvkZ+qPkCnQXEz0Tj3SW/oA+ayG0NPWM1
aZQlDuXgX1l5nQUPtVmkqWjvUbIHFBWPwYJKz3ugPdSiRoWO6PbkLVxhhjX2EiryqDGzlUn2p4vk
hFBewFteTZVnp7tNysacpad8cKUc5P6uHJ9bz2jU4mTKwXX4qHrci4RqcxB51mrlRPdt+DEjzHor
/5B9prjH1nzQhUvIrpQqf8qG9IEwfaOu5faCGYh1+r4oBN1kxrLmdOdRBpyC/d1NWn4YmwwWhL/3
z2d+HWHLMX52X2Gr7K8ksFrxD+FFEzKv+d7ubxCCPk+valwfnQsq7vMRi50Inr4lKiyEgAj4M7nV
eHQ+zjZpd41lP5kijHK64WsPRQq9RD1Z7Rqiz2nVnt53Xwz6pMg7AeB+66geUKga7lJxYtJozHo5
Hbu0GQJvukDOlcozUbHzpbRRsntDE+Xq0iM6mu75QCYU0rw6OJiVy5OxtmuwJGU2bTx3solyoKda
//CpFhtkEGIUKYofGJ+8Fl4VJq108OkNLlg+1IbRLuXyBqR01CT5kUJe5SVWUVFgZkx+vwrvpcxX
0IlhjVX9gOu6Rc0IQF4HB+K0oWF5m87yVOMbALeOphYABbR09I0DLAYY1yTIdZZYIsui/snM/OMA
/wvc0GPFiFeOnxV/95PvSRapH68keAIJXyTGXN5NiBMjtwWx/UhcEWOOtwwxFzsbsaA8Deuzdf+Q
IRn983/o9sBpaif+pK6CJk6H4ugCbjsTo2zVXJjwxMsWUiaHi4sUJw5FRwypydXGRg8sPHsWgu9v
/BRgZqb7sn14jd/zdjsFONKgjtb2dc1gV8rP/0gU13vJcm4ayF4YriOj8e5KBCXOiOX8kdSTjkiP
/rSbwutBGXmDx7q+BU6Fob0pqT/AdJH3c13OIKV3q9395PviN8a2bxkGMfXgQbkDxwQTLvteBvWH
D0+BjpebCpPiSPTO9E1hBi42bwdjd+1Com9PnV51fX25Cj4fPNBZ2jYrM/N0tfuvyzjXo04RVocl
9hUFkAe96AeDaX1VoZW/JkbHQZo6UGD0W/pVW7uOS8jJNVCWQpQ6vSHfd2U3jJhQ2jDh83nacaCd
jWcUGVk/poPUFy/t/ZZlu1thB8pfuEYTBifHf7244CMKCUoQXLqXqr7xwwVf50YgS1RdAwJWXAZ7
VuUiiG/MfQ/ErB9Yoq64LPxd3YxQKHAQHsljVBrk1dkYlQtukgCUBuxCpmLUQlzhoCCYSABpbBDq
pctWBjYvMIELdT7Bu1P361qBo5RQJ/JflbNyVEjSk353OS7u9NBUkEJnq9FcnCLLEiItf6TSrqDS
jW6OGTNopbIVU6Aq1hzhsHtFnyD4ittD/YT/NYJTsZHqyC4WllGGMjpayQfCmMqPI80iBwjmBItQ
WlTJlOJ6nml5B2xvRhD0/OxM4WifH+0zatUnmfPdZd4yOhUM7EzdwPKdTL4D2ocGg69NJXOTEKLA
KsYXfjRKSO2jBadhWLYK8yO6aSlQNyGOznUQyFNWUMAV8TRQ1fefue/dx62CJPLUebVQiRhh2vOI
iuX5iagR4kER/gY+3/5Ca2Bn7Ozy7KRKD98xYt6DDqOKqlysjz98dA54UYayCJ64D5L+75nncLqc
tlg7Rti4W+y0NMmx8dgCMYpzQj4mN12cuUhBWomPHuftwBmIlqMHb2ugyr1XTk8EekAS5D7z9pYr
1/yrU0D1TNwSYOQmE4oUG+nP8njHfnRwt0r7UP+Y+UelZtv51kLwovgHvGWJz7G2s7q1NE/+GUjw
/S00lvqeeisqFuS9HhrEiIR1ik6ZK/PfQGzzk7xO+gnbBdLysAGM+jX60JTa467qlTD2Z2eTYKUw
4wnRNvgA/UNtyiE/+wx++lpGek2NCDmEDIL3JUN2mxNE1peaOnV2GnnmQ7zGyRlQFBeU4wrFHDI3
VfSISaUMwmfSmGKj5wPPKDmWj+7d4LfkCpCAoIPi5ygftRvGkGq3OEQjBBKwiPah+VPpOgtUfOhE
aU7YAsUtoazNe6hAwT5i9ILpwb7n1xHDasDllzMIl1P5yPldlTF2yQf2xww66UmWyr/J8bD3JyE3
UUY8mTzB/ZjnI4zezTPGQQoS2MC7i2ywR4gqDi8XnkbD/4AuwVFlrrXBP+HRS25CntB4k7AE9Eu9
539D8YJPOWzd8zOXZwXoCZr07sobrpSa6lYHa7hMU9wKsgA3mbaWFApQulM4aytudPQ0+L5ms4/3
MxN4dhBkmXb0P8rLBOyGFkc54+E+HIi2GQK/QhXqG1GWFlY5ZcQtnWew0xg0r3522Amaul0Oityo
yLSXkCra4va13q3m+AIHv81sNE5ukbtkkU52MT8pJUP08RuSPNSrDAG2Kw2IMFIzsyJ1aEiTQL9Y
wFrF2rGlGjdKW3Py/OVzClQtxm1vvvI7vMqrj45FMP1iTT1rhoZoy6l5LRV2OpEHPaAZquMrgKtJ
at88SLrEYqbUAJfMbs2215gIRFY0pdL7qleBQop8SbWnmISCpidNp04+q/IjFU4jBgVQeYsbjgcG
wJxCQ9UG/9k5mksjvS2NEoCRHErYHmyX2kHyWkWqOlfOwD5VXytTYqGH1TyjOIBP5H2kvmQuVOkz
N6uplg+GkfixIIqm+iA1dX+XSAAFG1sx8rwALaepkpTaLTNS6Xq9c4EE954l+LtHuDoIxcQcw/+X
a0rUtvxsMQLG2/KgqWOhMzIeYT2zstlgGDJC5VK0432fP82rTaf0Ax8RxQl4vhT+LqyxeveIlBdr
U+wS5Kl7S7PkA8acJm7l6fq/UJsU/Fq9XeICMef9IhVn0eUCmUruLRv+GuQB2COgYXq5jsPZZ2rW
7N84lyNqqZxt5LfhnYMExkD2Pa07peOL42jZWDERboDGdJvNGJHIBSgZc9KbNZjihTS5ZvrCnKTP
Ay6ZderZM2yGTnRcSOSw10DdaH6D9qMklXdVGbOheBuPkF7GMHpvrfi5jPdV0HUFsXyKR3sTaVnJ
gWvyFR/1vBih52xDezdhxHYsUPna8UDclWDHQaaIzuQ7LRCL6c45GHtT/T2lde1hx1VlKdSotMrn
Haa3R26QSaog917wT50WGLOWLGmv2c4SvxLZP/0JnCnkKLitELPUoyZ2GtesnLbKGR85mtT504ge
5wH5N7bYF+nE/oMgmiC+zR+Kd0CK2p4CJIIa4yDLWF60yEA7UB4/eJOCjMNSssaay2RyXQtYT/Mi
jaMOFw+k7mVk/JSbRlST1GR/2GVK2L2VMcC5n1linrM0obrJYxSqUMU79jBx8k7sIcuTARydZfAF
quMyRBOKkSAH5gYSD65WNPv9nZyKJeYvojMRdFEgb9DNSlcysHEpkFp3YCkn5ltBD/CF8WfnNgue
DpnUCbTUWbNoX6+4S6wiuHJ6xu56kC7hN4+2YDdfpVAv7f/xmXPDcHJZlNoDj1kePfDu0KLVa+5C
iyLpmK8DR1tgKaHEu/tfkMrDfj2tKmMIWfU067l4eyy0CafkFQGOSabD+Sy/4IgZyJorcXjizljT
c5kTqvkJt0RsEJEWprkaPu7KJJ7pQv4HTDwCRxM6vHeCGUhmmpDGnJGnnueu9VA9EJhTe1m8alN/
4WJmMB7rnzIpq3x+KLLL/Km+wVO9Q9+p8cTvkFgKSHOXT8V/BB7jozBB69CeQSpXuiGv5PEMbOKV
cZZI1vrpwi+7LzC/g+AMMlidWGHSHCTIBOlwo3jzeDphE/kJ+MfJQHhkcPCBHO6Yv9SjMHp3BqJL
73F8XJrJQLFlYUh+kmAP17fvTyXABPF+9N8Xk9+QraCCwMMkC+MAs2d58hy/Y0i++bctJkv/Mo0x
rzcdvdaOMjw2UX3zANQAZzmHM7E30NWftLzQWj76sP301a8aDKAQ/LHUD1HwysBmFOZbKQSTwsLf
I/LNPUjUw7/XqPAjNASJ7tHg63YrNk6bHh57nKUgWC2JFC5emkjmVY+/7LX5AeqgG3npE1l7l3oh
KzIYslrw871O871MWNW+MXNZGCcGPT3VhoYc48dm8B7ZwSheNWywNJRXaRkV3O3+uSFTB9NQY5a+
jkqVhq6IrGWikHO4/tNBSr45Um3Vz7isYGzje3nBEt/R/J3eYRcuSEm+ZkPdQzd6e3yndgCrde+J
cYb+9KK8FVUl4nb3ze6o9PFKhsEnWnknewWjDymKfGl6UhNaQy5emiF40Jprb84hQW+ce8SJLOBG
+eRDJiIQRFRIHEPjdR12oYWbLCZqisVD02sGv2NPuC/ol7lWXap0YTELiy0WzYZ2+D8aGhMeHhpn
f83q0UIWaGAUVm4+rAudCWL7XCCFQlnxwcauiVlhwwfA4FL4+12ZhSis0kl2Y3ACi6O4DqBUQSSM
RERgItaOdvsTu2u15TipR1hVOvwhy45mSkfr7fbzAqxR9U1lW/zzzrJj7tJaN6Zb6rv+6GxH7N+g
alej8jY3662ChLClMlrIoZox2MI60fLP2kK9FBcCaDSI8L/S4ggcyjsUb+i3kT3kfcFttQDwdrPh
/AIHuPbN9LasG322wBip2BTMTcZrY4TmV10AcxiUDJ03/BBdIF7dgRUB7M0ThZiQ/G+a1w5P5cve
ERMzbMBiR2LVkkxyRCWkOuG80btwragxHDpeq2XIJqn+tAjiRlKgtl4b7ZJsYI5iHfM6LHHULa23
DS6m5v0x9vm9S+U/5di1uMvsOYbl+AHZXbIEc4nv6pOtgjns8/V1C2gH7jGcO1e2sQMCPrhajql6
exnhuxHsrDrVWhwqikZWyaVqaRSJ0ylkUND7HwKG0kfTq/uWaTO11IaN9gicld1yntjAJL7G+t80
RqBH6trtGl1PT3nVHZGgOj+Y4R0vxZK3eIPeJY2Utkaehie/LwKAfDCKFegMis49kLYS9R/U+68D
OimyUnkmZzRU0PbI8hGJmdUb4sNEV/YMbOBXskduCoqw8rxKTyudrR/3Mocp9dYuLEGS8TVRawbd
qAOIRA/yLW/u59SID4pDSv6w6HX2UsIAN+DejLwMFzAqU+zre59uK1h2Vc+J4vjywdB6QQZaItnf
5az1vfCtyQbdjeJ/qaHG6cKKkNKD0mvYwHSo6GhCtaY9SNB+3tuT7WTvGOqgZtOR9JHxbWKk3ByX
CnmdkaXwofk/nLRL7aXqCDPcyVSDMwP3jGhuDTmtBfpsto8EsuI/8sn2VXDVQoFTPM45h6+/Qfkd
MIHOI4dly7dKHJLALstKRFAejyMBX4g8YMV/1xqBhlKCEWN7XNRvoeq9BKnclcLBgIhWtqUwuLBt
vYdviAPTfGG/vzW6x1xB6WhXPP2YzxXQhZM5IWiNtDjvVlQnTpKwCrIIefk+ZXrkU46zVpEXFp2j
hIrCZPb3p9VkfsXnHhxdcf3/Ul2o1DVz9UyYgwR1qEQ4Z46nBuDo2QBCNFOYN1BZIovF3LptxjOZ
S4kn/yES2QtmtGfFmE4jm3v+htWMwVSooI/ZhuBf6qReATcpyIDqaHPGKb7jQrP37CcVvZWxCGRs
+BXY+/8tSNz5i6Ndb3out2mO9kmCwxwJTFfMtRvwDEmBps9Xl60OLlEx5m4OxaMSajCbYZIbPuYF
lP7ngjPNz2TjPR/lXRjKR1Ik59GtG5vbdWDoJFgTbbgQ6iHGAlLrVoL5ITXWdLFCYHiO3jzHKG/B
QiVrzFkFG1EftODUf8dmaLTBs9cJ4GmifWv3+kBbVxdhxjFB0I8z3gTe3xnKHqd2TkadyIWCG973
lpU5E5uL+pPOTNrpg9dbfnfsHLNPoq1UEo96pf6NxFHGrFfMSuQCac8mVYzggeMx9CwTPOYkXbzZ
KjXzcX0W6o7ygULomfPO1w2Fn5OCPRtrgQhUOapEPXga6TqqIH7tQeW1Slcsk03SPfkG01Akc4Iv
SuFzs9046TRKGYf1harLNN8si+lyR+dBJfvddF5JM57GqXikFfk6M8gFyRW/VVFKPKx66/KihkbW
oMeB2M2LSPLstnYZClA7A8J8mB+MYcACXc5F+wOENdHZsGyD9mPQP+QLB8ew8p5GhdpjirCaQKNr
99tQ12d0D9ET9uAXIWvwxb3bmf/L1ZHeN3iUbL3mn/3UWJDVvzr0GmLuILx6rYakre9hotbWuGAi
RJsqER9z/Yan9lld9L5ow/QHA1drMx2M4cMzi/nvUV4znEhU7q4U6mtG703oxlUZPnGxk/sUUbej
MERK1RGnVCPXbqHw4S1Fk7v6KurmqIEwLIyhlcfB6nGtOGwTOPfVPpZQkTrQyvgovlxQ0BZLYzYR
+XfEvwUTETP3dC4QWu1NGAqbyIl22FrGh3DkCLv2uMFb7pGFTheZJkkD7pmTbzkWgwkdsp+MbPlg
emRkOk/p6Wy44b+sh2WszkgS58zW5EJqnKDp3yA1W300vTFO08G38DmoTcamOpBREFFigsmHpHnZ
NG9Aw0ULGv1Gb0ZC3uIuiOIrA5fIe0mCZ2lfCVN7g4t11DE8cdztA52RWpQpSDClf9TDm+6Q1JL2
/N0l5XWj73VURDgl5d+/7aXfCBElxzwqL7ZHWw+lfdmzVJAGSuCQ4vf7ufXI87zy/ud3SRAEOTlp
4A/U2OdzIIoXLE8cIzon+dyl9l4JOnDPXxMreWwjKGAG0OPRMHf1ipikpZX2frIhPWZbivzjKKUs
VKWIOrnqe9+VYnYXko4QavRDA2jml25LYF/o2BuARtIW/YIC61MV9++Up50CwnPNYkupUxF5wapm
J4w+R5wN98bu/GDPjjQ+bvLdq/pDQjIYHVnfrKAma0zKWMiQHDgAQzWjR+d07AqYva2v63UGeM5/
H4/xSQzMMKT0kcmdOaVAjw4Xa7quRekyj5qfNXD9o+72+RNpX2/RuNyyXlN8K2aT6GdPFRWnc8uY
HuJ9IBZcaSkjKhxcXY5Hvo6D0ez0CGqfKjH4vjnS8XvPIrkjI4emcaohC+EH5FOjA5h/ktMKkSso
Ew1LPHI8yOUGwR1E7ORiwj/M9iPgSbopSGBbnxozDw+2nUEZNSL9ysv1vmHhkOtipHchJLngH2CR
BL905jY3qzpyHltRciuNui6cK8qULLsZrAH42zPV1osPxvsw2oHyC+Qb59bN7jLnOM7/oFiIf6mr
X8h9eggUCwHokf9PbDN1vsVcWUU6yJy7/JfmfmWz7A6MAoxNw6ojB6Yl4AN6MHHD3UxSy0syislI
1ya7vbjnRIxgFEQuTaN+3HSKM5pLWOu5upRkZfs6IN9ZE2j5Q6pE0kFkNYaOiB/E3L4+u/Jg1B3Y
uFCAFNj/Gs1YvOpLj/GdTR06YpVTiBBq3Hw2NTlSWX0PIQUFs7DFwDzC5wa3uKHB3XDtPp2j+CdT
JzS8UXclB8PRWFl3MTrG0ygPR6cVpfn/+8KViMwGvOw2Oz3xHY4EJmQh+Yzsw+AEqjB9ixnwXatE
aa4sLT2AYCBweLPbSdsMoZnO29712H218OrIwVVoVNaqOJTdFXj9XFND/ClsM0HhX1KB/EYKpV2g
s4KmWH6jQ8+b1saApfH+yyOd307DKdwGfRFUfhzdvXOwHDsjEkWRv9J9CrozUXWA7ZyIKOXXKwsU
AD7xSGrMa/I/Vq2o1agur669ucLb3edp/ftn7VuogR1c8lr0waQoKtxiqGYlno/Glnzsabpx806T
rBjk2zlYbtVBMcwOXePH98J6G+XUQr6t2CyTGODZYG6NbWOKcY5aXiTLeNs5wmUc3NbZVJY6sME6
QtsvboimgnG8BKyfRHHVzcxtr4/lJQsH53NdrJE7v9ltvszbY6ZCXmxRRz7+XHvh3VC56tOA9/+u
oyAwG5/rIx02vhB2yHEqQ0NyyXgxTSXw7Ut7i2giHFbY2d5QfRH6d86694d+UIROhb2CKegi3PCc
tImtX84VSQbpKv5I/q7mbnIFW5crS28ZHrRbzFm9ZBMrSfAYiTsowlwGnz4pVV0TlXXCt6dLwdYy
YFvT8LlvGJp0FrEDgVONl6OCt6VouiFKlgRzAd0hCcvPaVRVRBxzVOJszU9tAOY6Zzh0VeDkbJ3e
51oFA6QG/4p31o9Axz2L4+xj7vGW6vs9iWI3n25J04njJrfBUB56fylbtuUhtOpdKGJ4eTWWSccj
R0TXsaCXTICH14fqBSbqQGplC91Qe7ctj1l+uMoysl0UTY71kPVE+tJMCCZLJENbeqGI5W08GuuZ
+ok3QY1lqnr8Q06zSAOBHdsRJgQiHR7f99X+RTFSEh8RGMdI+Kh6tXe4zBi5PKMPrqOURbsIR9YD
2Bg+QgH/+OqWPXxhdzG8pA+ka0A7mv3L/lB/pjgOo6TszDjothvfttZ6g9pZ2/glM+vqCflnVA+e
19DKoxYiTqIjlQrXyCXOpRxCTtp1DP49z1fyc1orTHfgpuwxHH6elKEIgYpxN6sHxxoY+Zxod4gg
7QFm8VrPzfqIQMF8Bcn81I5FdXP3XA9F7WQbQVfg3Db67zSuoyxYSixKDi7V6NsqaW1PzonYSPs9
SAgaMt1K9osAOSEv6qDzsYwYjp1+CdwMWi2iy0F73ngRUwbjWI6ccEuJBEHG2PGnzklec2oR7Nhp
XTtAHDQC1s+LvCaUfcZaRi5s9WBfI9ASsc29JLoBHJI2ofpBAa5tCdfQhOQl7OYQkKsFXcnHiCJ1
QPW1e64PPuI3Tjgr36cOCGNDJo1B2L716kjfrcErOvl2gdEA3TD4D2P1JfmU8da5QorSc0KDhjYe
fR/fnykXOE+F3D5C2F3sKMSQ3moyGs0NVi+79AJFL9Bd6K51ZFRI+QXeAskHWmHlziEtkDBeU17+
SHcZtLUpAfWvtF+QR5wlyk+ixzD+qXAVoU0AcmooFAPJzrwO2Hhfudm2rY3UJqYfaOgvOCKeSwSm
fRPEhfO9kYgnlEDkZlDMfNlGWntoOEiFKdefzIZF/qfHWOaLVhVSATZZN4IRhqJjxj9ewEa+rNr1
kUjvPZzpgfSDbqjLn07JWKsRRE4Oax/rNaWrwXIk/F2wl+bBdZ4eTwea1iGVuB3SqKuwTNgWnBqp
9Q0YLO9cuzYFkKAr/n1vwnXVfFaMwXjhw4EViBe7Fdqkl5RcThhfnyb1Tx4GH2ASebP10mIx6yNn
oj3B54W3/pDDXgDYaydcQdAOIieikPUyxYjll9J0JfuGUzGpXonjvFqBp0XEaOYn6/M4H7/3kVK0
Nzv48NCAo8xlUkwrTTpHnlDsAHjnNQoAO5qdNpTBw26nB6JjFSKlnU8Ton8t8kJNWpBMX2nCBoFU
NCKO9exW1g5HDXSAPzVQmxJGuuDpGrHPku9tGiargK+vjyV7V0GSUMz+DqP+0pEBhjlUVWbCkgRg
KRjUrc43FHJmVwNfvLwPyfk8RtayQ1uq7Ob9GbZtEKQeqqYNQn5KpWUqJfAVH+tx2RIMgJ4xaOLA
LRQl0tWhcElTCYELjFgFUebUAQjwavuX97y3t59OH/2qZmnFb2XjsRlrrfQsCNr4OlRVQDsdt1P5
W8v2DJ8kLGgqX+qxGan3OlEzHsHWUet2ssYCC3JID6QGqCwlOicLiVP//sc9YcN5XPEPZKAvaWv0
+3UUeMIMoQzADXkvUCc3bwXCqsjq0pCUgC8YmJZ4Xll2mhCMCMGozu/k92CHt8W78JgkE+uj+f/O
XRZlvmk/o3NeQRnszycV6IyWUXmy+Uisgdmvb8Z1FGyZQlsmrT9kc+YMsy9DTmz6hR4HT6w6C5NE
9SflzKf+tGeCESB61eGkKJDgqZ9MmIJLHmFe7Q7kPQqcip/YHU9QfiI9uOXa71hWA6fS/gBEvKsj
9bdj6LyjY+NRtDsiXPgbHZRTyXuoz9fMmHsRW6eoS5zkWkLWkjDv55LyVNAZz5I5YHM3o0zpxNMI
BMqvyOHr9pkHariVX/7aBwmKTwej+CbbMcamm1WYTMKVy5eypb0uiF/rXxE5y3vgEcF4sQyunXAS
j+zmEv8fff20tZbzYrO0wDjp/p72K9yzlPeVcD/Xjuy1oWxMn8FI9Kw7ggSJRz/RvcSMwbWDdIwh
KDMsK4Ijx0Ifa2SBIsyEP+DEzN9G6tLTdDA/XPhlGHoN7e2n16SDTVUILVS6zoJQs2/DCJRqScLx
yYpqGbfKtnsSEAqpJBpQuoiRcmxo3+8/CssyTlHBBPMT2MU9e+Jtv8X+pxpf7ThtFPrWY3dn6MFS
wuxw1HDTI2x2ICd+eg+CDe1MRkpEYma18JaGDsqXdnaWjKLs2CU4lq2b8m9HKywMHBQSSuD+A90r
p5C0FV2D0n79rk/z3IjrqtYAe9Ya+6k3uo6JRKth1ZZKZtk0AntX9VPfWfxEHEsncG6Tn9yjkZR+
PRCfa4HDgWN1dutsUt8bB4K46/oKK3xTy7/hGsjbwOzESy97xKmmu5ix+trUcxcj7cOzAAiowCe1
f70wJpfYDAA7QKhXfqMvcHM5UQHKz+0wUvxBO6m66OAABDhkaKV9CUNLq0zmQByIOThq2oGJyGZX
IIgHCpiKGo09YafB630T4snLLNFsDVfMMxJZb61zsLTb+lBAXXBsoBNi/MZ+ndhvla40S3VMGcoS
yTPEIc9ypSq+91TVSbhwZycOdwUq+oCCvB2pjnTM3FwYROYQFMZVZ+UXYa6n+HXlidvnNAA40AAC
nn9/3kBluAfbCp8QD9E1Ir6OKJ3LKHKo42A9Ixdjpx0dNTmX0+vv5/UirSSk71LATYY7en15SAcb
/7eu/pGAIFl2AqHYraOTxoMwijqpsRPS5Xa65TIK/ooVqJoR8YopdLAoG2cMohTy+yykJVbpgu5F
yjhP1D2em9FFeiNjiXVYiaB3uLWF0uDLHyRGesy15tPLVEBiq1+C92H0gZWnzgEGTu5AgSkoA3SO
7NnsrkYEYrF5iRMbBDmPA+58DkwUwYGTLxSYAqJdls7/3bs2w/djNuS1SjTPv/c7p4o5qOaUbenr
yonvUMA3626QItmKjcRKTBt/k7fqzax3cxAjQQnpwfFidQF56SZXOEEmCUhEp72vXpGpgxOKxY1N
VIrHonqDFjSNOY2BLcQmpfMs6Xz08kH5meK2gTmzHCRp/xQSgVst6xyJ7lpLCN0sJBe0t6aNEFCg
TtIH19qk9L2buIKlB4oPh05KrL6MtJeIQzye47D1pVJCFe2cHeWEfQqvpsjtWdvpXeveX/yIULV9
hKqM3XaBE5pRGwvKNdYpoyGxHHldQRQFYQnqcczPK9n3tDZlXr/7QCPIOnxx4Su726Qkxl+WxP7g
+2hIe+eFPYci098Buid8e1ScDsI7X7kqRVSXexFpkZgIi4QqUN4ev+LtkJh1t4iyuvT+wS8u/rEu
BTB5P0mtKG4616mKRvTQIloHvVMchIeSSnwVLBTIMf9sOpOQUJCUun5FQbyoDDp59f22yP53W+SN
zYyv/sK2CM1Kvl275XlHvJj0bWbfkCzWGdzYji2EqWYMHXoiqDi4IYKmdaL8ZcmP1MWCmyUMkehJ
Jx5QxmdE+Db7pMYmDx6LWb0QtiVnCZm+sJ7eIx5SecK+OEEqcqqVpPeDiF9ESgqjOUfNJN944aXF
qBzySQdFea33e0C6NXNG+mfW+Wut8sXbn8blWmbA1d2O8nl9E5vEucbElFFnoYZm9u2na0wovjE9
wcUb1ZVK59LASxplD/KTw3+S8V2OLHbwuQO7KwpY4V0UnL0WCe2mSHrAR/NnH7ThfwzwQToxq5f9
7lFQ8/GzdbQJImY7E2THfUaUnuVnOEEHc88345t/7WUyk9ks293vj5eT+UsfAP09wKJZDTuzGRyT
9YqqPRTfairhj8Ai0coRKV63sOgMXfAZFdYuR30EkjSLT3PG0W5gQ6aLI+ejhxrlreaPWF8aatOY
kIwwQKTEmDnLkTk9FN2psOAT3nRvnBUz9gT8EjCdMXm6kIRxPpZ9C2nCbme9SX4YOAovRijaLxdD
XESb2DSNggIBXkUcHpmRTnH0mwzpjQiTBoHrUOpKgDLthy+SsvLOexANkshmtLCdCoRjZ29dBXcC
BsPatSZpDMud9UwN1x3qmWHCyWWoEUNwKiV4re60MOGZmrDMtvd9TeoT27NEu4zAzpHTN62DG9ze
Pz19V57gIzpqORT/pYdmRrYrvbzghUMAhqy6zUJVSnzU+4haiZUB6C4DtAjnaaKfXdYzPYA4wcCv
K7v28H2qQC/JkT5buA5KS76Y+qfLPm4yZQyTzMtJqU97il0XLOsTM0s9KZVetMbtCuLOx0V4fbYf
g/6Ikv3MDYmXwk5IjrkGbyfQ84mWN+GMeQIouY71xLbum3k1Evwtq8iPZ/puXsEmBs+KBNvnylLM
u1KcsEnL5FtAhwEJv+myvZXiszeTU03UdNV4rQ/SUnUlnWYRLq4NeHEiEtifY63BNWUXKC7eF1Hq
AYQ7wgbtX1ipBwhMbTFMMbspytqxQM+r0Nkdfpbd/tbu/sKKc4/naLc/TqozgPQW9O2tdl7sL69v
BoB+UZbhTZafkNKit/rNGmJFvrLrY3YkmdxrZ98DMMu435o3gQoEdk14LgdaVsdEzHdwtRgscVZS
JEivhQfgP52j0OKQ154s+yucnK9P6CebASmVJYAFXJSBb5BQR4L+Hfjbyx2/ruuvvpwqW7GheVTH
bc6YdGQw3/WvKKCO+dJKO3GSlZhjlp44HnuuAVAkCgQnlQb1b7Zz3tkUgVBaTz0L1Ad8Vs2rrHdE
xJUQHw4IfU0cjBh37LiDWFAlkFsLoeejA3ckeYkWTvn2jzfekgFnLrrqgggITMaYKNUCTJ+KzK3A
yTVEgAdhqtUhfsbrJWocI+1WGqr26GKyUJag3/WGq7XSxFpFGrxIuLKzuPiLxe3rqAO1crDoHD8Y
Ljj7zSqOWUT0Ly0rNN7/xW7HppP/DP4JVeKIKRxTZHaJkVj133uWu4atDFb2GrnJhOED8FL/4KZ7
cTr5KQlw4LLGdY+RBv6RctVGe4n4QFhDmMqAgBbOmsRGI/hm8kF0vJmmeAplEoxPbL8UYT7D6YFX
QYesrCKQr+u4eLhFA2EPkzdNJpyN4pmMqf08XTicHgCagQI/+xRx8vNFRWXQxmiFztzu6mwh2KOv
Il7smMIMKGPKlO2OP9x68nBKfnHkKdN+f8KZWNZzyHiiUUjr4auZpNRRzS/Fse7c7NvHUavsZr+A
lJPuyD0BScxaUtbEj3d6kWLW6aMgnkN/OEdaymUA4JsEYIziogUk0hnjTX925s4sOIF+YcKU2sir
3QzENM3bjszYWuqaV1nGI9XdTdpUbb0kCwOLVmzFkG5fsk2QGgYoPab4SLBET2p1xiOdRzNXLIk6
XAEkpzCcnYEfNOtb0YYnnMTAVhy9VBKmErcnBs9gPZVI6QdFxijcW6ANiquFA5f0BMb4V1Byo8cU
ILCUTiaCkC7YWBoUq1GH2wV8fT+wMI1wiJpfCqAnOhSy1Yy9VLKTHRiCKk+xSh/t6KZqHGNYMBk7
rlOsFmXLiZwvEwJINhO4MlU/i1Tb4f4TwADcuiHHJQTpiqcdgaSE/fq2VInLR/LzHhxIR4uTvHp9
X1eyjB1Ez13lnEYJXrSWPspoMxpEhJx8rK6ulZzuyvRhbRFmPGq3jI2nYACcaXc3GpHb988Z0fkr
bVVTC/WEN0ezZNd/KwEaxu9hAOgSWurZNfmVi7SIEw8KK/ONo4BLBTikSilzU1/+Xn7IqJjbLkEh
LATKCw9jOx2elNO4Z1zccrry3wTmV2Sc4F3ToeLiyAphsI/b/cz/NivuiytB3QX+RPr1tn8p9Yk9
VS6WdpbX3VJYl/OytdYsp/y3u9i4CmraDxQNWhe5ldL4Rd5r6TYpKJd5K8cOTWsSa56n5iVT2xHG
UWXd0DNz9el8lw8bmYD13ziUqW9Qw7ymaQE7kozUFUYtlYlO2eP0uIs7UbZVcukqbIeGQt+lkiZK
ZBugDVvPg11mrjQYR09uHeogNjReiZ+q4u4kKA3UjgxlCK3SSpZlgth7hHgjq97SfuNYxaOKhvZa
x0vDxBW11E72NXJvjoe7Z7DlaWp2TvykqK2/Emr3gXRtNa5w5KbgKbSEc//vgezQsw7pyuv/+yyN
QzWBbnhl4mP3L0lOpzNa/qUfj4drEfCbbVAuWp76pYvbHiM3H4vqbdJ13phgoz1oiRhHk0MkBoUe
0xGyY5QxpVl/aepF1vGBxmkBwZ5X85/Gpciw/4R2BzPDrlpkp6ibFYr8nIAIDV3Tk/QParJ/8g4U
l0k2DaY/y7x3ODkXR+rjZjRG+dvcPbqUmwQdE8F20QaNCYpYt83tUTIa5yotM7O6unBoF9pGvRfp
OHeV8bD5J5qx4wFY0f8U3Q6rn/5g5kFF7vGCLSI6eILvZaEpbxCCRwNeo/TcUXt8ErhNewbdpOHf
3wDFu5Z5f7SVuCaaQBvIeYx5BDXoqVb7Z9xeFDOcJp8ArRNx3jOCzqQ7zQY7yWg5ObLlWX3hRK1c
Dw5ZN8JjMkLMaqggud1ajThGlFsN50s8dsczbrJYedBIDwQhTi/tVc1ZsTywDCmz+4q4nmZXLhvQ
HYWxOgEi+PWnBJlWnnCxe6iD365ffM4B3jRQ7t9DiJz/mXMOxyxeSOV1jmicZGfwzU+ZYhqurnn3
uYQUPt/ooFffdDRDX33lgKcZmr203YBNm7l/++iybhcGy8MVuWNTMu6lfPmHWdVNPRRIKcmjdmGD
TpbyUOsBWL5hBR7WzdDYw/DEKgIRWsxSn7hVXBU2J+Ywn/1gWPAA/YjS28TuuuTGc44uex0rIu3Q
jEbB6q1AjCW31Jh3u0d0eoSqvj7QcCg+Vs7Xs9O5oQhU3cYBaWwG+7cnw5gn2qjRxiDgLU8JEVDc
66LxhNUX11ES7xrmiRwyn/tDKMmcLdeur+6trSsb87b0qfLEki6XKxBRdITXOLyAR1+EuHxRZsuF
W5AWouzZU/WJ+vN2dpS5RZgOrk7HeK4w7GW44MoyR3Zb+ICuikJLRsrfzLiF1uk7Fey6l3UlqOf0
Yp/srJU8W9D2jdpyJNmI2TlF9MTp3LIlg1guQyUe0GZYJFdwzwbxOyW/8Ni8TDXl9aslUS7jqFrJ
6ghfa1I9CO0SLGUJKQHHibQtolq6PBl/TDvTw9mSszPzFmsoAxz7ZvQAp2aiphXqpLeyB6VTJrSa
WuUUqLSdwwoF8GnNVkugAxX15z2pXYYYndYTxhZ01FaZ2eDG64Fau0wcicmsqLt5LjMNCoBt0/uM
qjclzFb3aRW2Y2U5HPbOyfZYfC60VfVHqvmRmRSfIDOg9gqu9fM0WJRbfgaX2Z/UbAwYR1eZFr5n
y2mcJ+sbPy3h4p6RcCEkQMlewCbPWP897RVHY8y6XRHHrkTBxp9KbA5JE81vRzrLIWtrUtPlFVmv
5gA+8yaZ+bJvomCmmehOH0alBabmDPjs/zqVhRwG0kj+LVicwVzZMuvdp2W1N/ifRVQhMwWUpisz
3TYimRRQTpsGavA1xQfRoocD3jSF6Cw3snpDswQpCPnajeIq+Sa6u63C0QHbF3Ur7nhhDPZRFNWW
iCHONRAaBxEi3sjAixULbRXi/jPsJJJlXhZWb1mlKwCu3CcU8tQt+N4fj4birR0igrn1foq+3tOm
/UzNRYG7n+p5zlOA4Yd0HlXJg9dzO1RqrUQqSeKztT0byoJU0TPS7SyjOqoPV4p0gLGmN02FmUp9
I+uiUkh3lMc4LafLPzbzhsAYCU292888ZFslVCsteN1SNpEvwTwOKYjusn5iDmU2wKbHzBt9fl5m
ph1YMY1UD8cYgXqCBeBYaQzBkMSBrCQ2jpgA667VHcCqITHaPs0HxnxSq+aqcCeT7EUZ2fbiz1fm
3BnTXJ9qhIFPjcBBE7WTVncQQMT9kprmIJefhmbGXgjia4sK/jOAeeqs9ZLv0cLyqdDv2w3cki6g
/bm4aPCKwhISvacOEf+WXgwfuPHapQ80l0lmEvEthdjBi63iWpId1dEkoJyJOsrfmpo+nTA9EuTC
79nKbejezKqBej7nXLhZhdu2vieeMgoP6ULxX2NJajXKQT291TzpeCg6nyCaLoD2RqvRvWdmjZCu
nSXpar7yU9e3Uvdu41CueuqL0Utam3m6iYl+tBAU43WfIfBQWZbVpYRTAOfSe1OQg7XBaZ6YXpBQ
AbmH/YfEgk3BkGw0v6YUIIzBXMSWIHBzzzFr+P9Sub7vCIxTrvVMfWM6jySxUJJMoJrPyNQnfZnD
qZ7iSzKLuZsVI/kJKt6qC5kClcDXXZekX0r6nwjqnpPAc286DM679zC1VnS3LIAISwm/sEocIqNB
n5hnLWCjf0CXezkVQDguEB37EV57aNoaKnl6mH7NUuaVvco1nsrJcgu3iPySAtr7k70VcK4QBleK
GrqPMbQuGdl+y/jM2R9pgI5KMU3nSNSoGij0sPyLtLnFTy5CcxHyOXKMYliQWCpbCYGjHo5L/Dtk
dA2CJlh0d2CmSiEzM0MTPhZZ9XN5TvCH4Zy0jwBiko4vsEZpuhmg0dGMZUkGrHaMicFKhORXfgnr
YIeZuQlWdF5gTAmfZNyvyV2fjolWGDDV5ikBqct1Luu18r6f2PNTRVnQB17xMS0vB0ha4gsoZ9Pd
XUvH0zCe+qXK+Q/gVdamcwtD39vBVW09AA/zbXdpDum9GO7JFLF39NtR6mBNZrLBdP1XdbNbvXvs
1ueDpVAuAm9IpGWzMYdjgjwfyXPvGf7frux1AU5UtdbQmSTIGjbK7b5YAVGNh6eXPqwh+B2FoAiZ
2ipnng2i+lJTG65Ct4942PwQNTeMlRCbIVomBHm2h8v4RBeJUrJe/9fG6yUCPMomkp+St+C29AOp
yxY9jHn7Qd+6T7Dr/IdLlWHsyRkwKKFHvTSxBfF5q6G1N4qXHvpb/YHpvJYQxmtTHLgtGD0B3jg3
cOr+BrRim8oYFL2dcFUXXu1cWXjFTUwB1JvEz6OQqk6YZQJTDtBI64hM/HxTQ/S83WOSzcRNqVPf
vfpZCU0jrKpSGQ6WS7lR1JjH9ikxnAjBfNemGbGf8Nd7JNuGNtDJ/XDCALwclUvjIfBpapjz2ysg
8M0Zd3/Lq2Kt9TkNu3noIddYXoUdXX8lim5at4OPoJ3G14vORyZvpyiBjckEyk+CN6akHv+82yK9
pvIXw3bbpJWXoPU4FLmZ7si1pR/wbQZaLX9AaJmrZMOmuzHFVgXfsMinxzaXkMVoS3xnicOiXFId
fzdNP6MYU8gpe0NMG0T19IFyLGJ6sB5PlLoxXZsYwlYug7Mqwe0h6AMXiHV1xYseRZjxmUAwC1Pw
fZuR4iEK9z6p7c9JiDTBJv0NrAUI2NR4zz2yHhjVvvB9EWo0SUpxGg2EXfiuAfP7EaMeJrvZAhPQ
sWvZsNVU5r8VUEEUp5SEx8JC7bcw8s6ud5xOLYsd7wJzfRvXSruGXuGAHWPSVigkxU8+qbvStG3i
4T8z8UzvfQ0feYnlSIokI8itppA37DA1dlhqAucOjnv57YOP1qH9YH7ImRE+a5RvHFQtw4uKK4AD
yZ6YllLYQr9lZ97KptF0jPFjA3g+i6ROZxkjdL1UEyd+jWGPTgFg/4HnKKwtvlREEVsw0NM0fonk
1udAHuBLxr5e3Sre6351NlkIe77LtgLlLhg9uJimHiUTm3VJOPhPPmZ/Egj4vRo+Rtehm8QyTMLd
kgTzjS+VhnaC5sEQoCS6xz4VnBCnpKF/RdfoqJE7ADoyBCi0bvnnJ3AGfuB8etW2txnG11B9QZom
HFzud9GXMeTKbC8QoM8zcdgxfMrhrAwfEYcWeWgjUMATx/x8J36ZC7eE/s1DE4q9gs2tV6eZv+lM
z9BSXBXqKLpgVJgwfcX3iNtljQGfDuq8YQ0hx+rExujAhVkMT71xgZsj3q5wcQNyWNrRhJInk0wN
8dHjARHJf8kHDAPJ76Z3EHzS5pTa0ITFMqxyFxQJmcKGjKAE0khg3K07cSvYqMyPIWb4RCrc+5sP
8Aj+Ne5poKRbNMTCqX//yFo/jnYacRbHDOJr0Li32npbfmxurvwlCSfZWFwFrdHUZJ+PR2Yk2v9W
LqtEz+OsRsER3fmMC0yQuoo9uaq5fVUD6tBKs/jTa5GHH9NsG1ph/SLNLf89rFaJ4Uf4n75pxIrM
6XvzsmtQON6sMdQhZ+xrrKqX3qr5akrxGBHRDTB+jDprwyRcQD5qfzGIxGOsLKUJl1SoJn77DZAo
9wNmOsy4PeemJ9pYVUZhhGibNYWqGmFCFEbkJ9AE/qBhHhD3JCSHAJa1y0Pd6/g2Yqe8GsECoP7D
XeC1vTUzrCtIMxFez+Uf5WU0/doWxZJrxxRniRiTbxKVZUhBEw8vuw8bR3CWd6npWFOYbQP6hsxy
h7dcYzmZzargelj1hMxo4RpAFfsERrHLuJqbv7WG9QpMOmaNhgAw7rqR0vKH5GGboo3aCC7FEg5e
BaEQ/mY/RdtPvNR6FoK6I4ifnKm7yOiLElTmfEsWD3pVbiVH2l+Szlc4HVFaoRs61+RxKkdjRSSP
SR41bWm84+mWvBdNIfXTVNsaBNswAsliH/QTgvSBY3MmtpkAZMAXF9QpTks0R5iSCgtPcUzKviSC
Z93qI+fxJ66ROPKoWnW3LZaUwWg15xfBe8BZmScFEhxJzZ0diA5ZJhl9XHSJceTGLDVdqu+pjzri
FWvy83Th+YrFF4b3vU2KN6sct0Wh4TR6ZNcZlX1osmjUV+/ZNVC0MLmXjNStxB82wEsBfhjJJADa
fS8rzbIBCwcXb/3cPS7DXyM5drho+mUZHeDbcTrcE5hlJmsiybHRSd/GkmIHg4RkRDxBQRXGPfL8
05w0O7MwCETFTzAeQ+xjThZhCSZKa14dGvrWiurVI2dPr6uZZAvac43tEr8FHvhn8M6cDAOaeSqe
IucjQeOlIrQ7ow7hH7Fu/kn8wIfci+zLBogpm4QWg1dJF9hVflrRjAFDO71WsnKDrgCQfzjuVmRa
zXEsFd3xBo6bM0usUjWUHfxm3ehcGHBYFgYEEgHCVwIrIuYrFucRMuC/3xJEeD4XH7gZ6JorJTQt
5QNyh6a/DQoeFo30vs1YKlK6h0LtCGA7+jxkVB7TYtR3V0ZbL4I2HQe7r5vIfxOLNQ4xcP+yuwCc
lgnqKtNYl67WbdB9rJDOMu1SFr3dbYw3wMlXKQesIpkuYA/NHAQ6XFrdBYKi4BBN6uzHZOD7iWHt
7tTj0S/mb5OBckKh9WRxZ6NiMRmRqVUgfiVC3mhz12nmJkPoSJg8KtO81fQrljrHjwb0M3QNgWaM
8pN717XZeVfocKswKX8r7ejkpZlxE8nbouXsQ//fo0bJUT4Q6C+X8C/uF5/15kGrHm2HqaecpZ5Q
JntbZ+rymW6ZlfG+VdRP6OtIaNrm02evJQen61Ty+ZgJJspYVgXaYbUWpoWO7L4J92M4MRHLgZuU
pctkOTdGy4VJ7e4EY9QF44lQWvXbtcMDuGueO3cbJ24jikOyl/1sKjtK+nZkrHRmdl4HrLdeJifd
mv/VwmY9PsZPAGe2oZMhqJSUdsplK/yIdnURysgflGctBKckuHA2B6UmDTxPRmZ9WcscAjEM3Zdt
EXyq7VRZ977NC+qoVTznOor/aNiWNet0UcNIgmTVAsOaesV4j+ZCElfVOQsKZwx8u3gTNJHLNF0G
V0L9bKlGN7M3BTReLw34ouT8A5lSP6GD7YwRXetUjE+wj++eOP17bCNOkBeBhuoVKopLGc3dFiCQ
h/IfVzgK/iDKD97drwUJMpmSLGc2S8vo6JodV+3orWoe4muu+w4Td10ag6AJ/cHUDXPzKLslCyg3
wwRLOhXRCTTO0AF20omBUrrYqxVWWu0MJenjdB9skP1yH/x3TwAcQA3evgES4FabbZ2pjJO6RtyD
bvtxuC4ZCneQPfLMW5uNZR8qaZAR5awOwRhmyvjVWo6OdS+7DjMjj8H8yivkz5rD2QDG/HmG/xKS
UOIIlK+hVXtI2dI7lgbGav3G3w2mpTzOziEr/x3/mE7pFCnt8swwbMR2rladg0mmGi7STyqspeb5
3OxzZIvvniQFOU4Df621sXtAWRP9JDgi6BIilWoQ7EEDXlvtKwxeayGlXcaCcH6nGmT7i8/xin/O
BttJ1G6AyNECbItCSf8trg+j67UL38syU0mO6onMvYebRqu4cXpl352NsePVErfkA+8kv0SXMy9o
wEuHUq09RvgHoXioViwzgCnszaKMYMztt9Fml5ZM5eBxih74IlBrgs75yxV1BJ/LbupH7dxvNeZb
iQqh/rL/1YRhd9t4lU6eLRTrKoees37FZMbG4L/aoYvClsc8WfxnJrQ95AJgxAduOw7Po1N/toMj
Z8L8Bq2x96K8tHPLUDm1nGztBhoDxewvSeJVTPTeBdXfT76nOB5mK6ZAiyiHDLbMH+pPq3StkE3X
BVYUO5V63qgNlnr64nQSrCL2SGp9nSvliA3FDyN+s3jdteOx3QXp909Bws0ACzIGhgDNYgAl/Sr+
bC7jXayqx3uCjYpDIVk+HKqwdj5+vw2K0kVAWTO93HkL1TKLktxLiLOBqQ3S5aa5+WrklxNJ7FZG
+l+ZPmBP3pqDJ2vOo+hKKOdz8WEySpE/zHrjdfNRjMZxcMl/8OmzfgbGT/r/92u95qLXlP1lyvwY
A97xQp6xU94gq5xoBiatZU+OjtDshSVnZH0tg9BIAr9ZfiJK2PQHxZD65cBttS69KY+h7JsZQnHS
ATFsMvat6g5PYNw+/IDQyBxpEEAtvh9srXYFsyIZAihDkTZZiCYgQnuHp1IM8sLHSxuxPGjzMgci
nFxi5/NxtBiazEhOSvkLt+NfPQfLAJjzx6Ii+60wKEanaTXaOsZHRm16umEbkNfKKBFn2M7I7uXd
JP6mo4fSL1rSDNDnSXplChX4UZpmk8i/RQoYsp70hHTX+T6Pj/k8V7zw6N77iN58ohZvMkRD3WN2
0YK1S1wdqv5QXoqD/Y6fu/j7GDO499/eE4etUJFnBWiiS+DGRwiG+XfjjjhW6yErS+NWtztl7kiK
98MjLYRyeO5epMqrijwEKfrwQ8FKlKXjsKODXdmMhvrhUFosl1nrpgw9QvkbftRNeS2DIDS2ZH8G
HUPx28genswdnZWyYLpSi/aN9y3TTjbFJKA8FmI2FcTtD5VmQDq6JKvggKwoxr/bLSS9/4FQ9mRc
Ul6uDfZ25PbypdJCEjy7WT9Ai0VLmUdW/IbRulVbRtKnXcNdxqEqyPbGU7HHiguTn53x5aevScpo
C+/OgET0JLZpRXSTZ6vmGL4UtIBlYwwlOyydWemdZT9S9yApOcKiTp3eKvVdr0UJG7Zt1M3WyyEM
t4qMwzcFncel/OE74JWOsu8ef2aI42eeJpBMz8gQtxeNYDUBXHbSv9ZsFEaP+6PE7W1fbXaF+rHP
qtjB/bsYzfyFaKAgW2uK0xfWkayuCJ0A43zuVGiziuHqolpvSYty5hoMkDN/GdzBRtg4zgsPrCBz
dSGBtkuJ+6Oz13AB7+v9fYnFu5PjRH907PgLJTiMrJFKvpvg+XKjQNNVc83lIJ9T4F7JuKmf2Tn0
vzV3DT4RKhQcaHW1ZXUA/ehraWNW+qNvaKGmh8MqTupftTK+uGlz8SKYeQUo6HEW9ZgCeN1CVY/p
015AnLOdJAeIY0M9XCVoTTWUMElSUBPB8TKJskR9PWk11sLbqkn89uJF1QJUkG2tlleHNX/EJMWw
xjWcJP2B2k3dxG5LXPqaP2g23ULbmp9ROlTE6y5tcn5olx/RRilxP0cSPSaABIlt5RzYaX56lrkb
MUmHE57Dt3z9mcFvLPRzgVE7culw78mN6qVMa20CgGAC1deCiOE0kNv9VHEemKwVk/lmh1Meal3f
bfYTDGzlqNX3Jkiy6EickpFTfvx0XMy+dcoy9XD2Vvyrj/S/LSrDvsI5lxM7v8Uz+gyu2TGVb2TU
e1mj92jTv0vX2Bsk2GvK3Pv8R3JPcRRdATbyotcwnJpo6GemZOTJ4LxKXxRJ7w0MrJRig2YSUz9j
gFZdq9ao1zSGacRWQYbUX60PJDmsPO/8P4OXu8O+7YILP0ob/nlAnAJj5C8srDlWEzYivTmfrbqC
2K3fxLFF6FKYibJC6goqjl+uNp/j3LwuMNjqVWhAzGP7naprfZSrT6X5GM9tMJesGGe+6YtKpZRG
K5uAw8t/txXlRxv3L/GbFn9fMzlJA9E5VoQ8RPPz4u/8GDili535kX+SMSbOj/6UBdzWDKYAnzeb
4E77cxvPbQX/ZDHgZ612MsZfKlNqWKSsSYmfrX36FJbp1vTNg9bRWd80fFNa9I5yveKAWgh3yAB6
8o/w4Km5e+t26QYj3xhqI2yjw8xPdcdVW4VEKy06oPmrfJdsuAQbRijrnB5YTw4hXxQZ9ddcDa6+
X+2yHrGUpLQCDrTNeuqZl9EkPTjCMlu2dESjHlR+j5VGmpuJxHBdNmGkUyKdbzkqjGx42gSbi9qV
j2dZLhLLxUAm0kP47kXy9rld4lxZ01jlIm7SRXjkkeJN1RGwSoyGFJw4z+VgvCb0hvM+uU2IZx0U
gjPjImjQDWhM7N2iomMl9NGrXIcRR54jsUjm8hPnS1n5DewSzZ0c5pHT4QMrvP7nOc7N9Rw6SZQN
JECwXkpBR0M80ColZ5fUWeN32nWbsETwBXUWqO22lru9JftV6GzQmUde7gzgB9NxaK9p9knmLhWV
vGUWjR9Hx1ZHX/q0CRpYAG6m1h6LBH6X1zn43fbVjsgYmOWQavXpkL3ungqKFxmHnFw8UbCGAI6v
R0JMjHn3huv1FdpPk2Wur2wyP8KIT2D3uJOXS64OPP1crksjiFmSnP0jISKFvMdu0yaq8ouPSVt4
sWobf8AphVDQCRmOCiyrY7+94QTlX9/JesJtxGNjrdbKTxFz2z90zqswj2z13c6yvWSw3dsEy0Gg
HjCU5gQ+1PgHl1GCv14eKm9w57yCo6+CWC2UHB8G6OFG0Vfcd5c1Ri1JrdiX51fzUGfOxn1lDN1X
T8YERzGFCb9mtv+BySAZDY8T1LHTskB4CsTve/TEB28ocJrV7O8Z1SHV1c8lepJIz/no0QDFk3uu
3qg2Sdyi8+oo18zTpAYtK/MJY/mMzh5Kh3ROd/PEqWxjzAr8iCwNwtmToNtnWsbhYGJSAKLo+PTK
zvHGd1jvCVatsh83+kPjPUxZ9zi/Q/SDH0/hjTgmOzoeWp1aZpYk6Ot0Sbx9Bnz6N/rMDG7D8GSJ
9v++TH7lfEz6Mwi3ojuvaDgu7+vBcVvV+BzzDNklFYCbjP9Dq3naSbdMjUD/FHRvi2LTspBEYJVy
7VMU0ebSbc6zk/0gxKzSoAk8zGkAe6jsO9mBN9lvJVNztk2kxp2s+vFkUViKuks0mTTQnfPr9SK8
xY7RQiL9tKFEYYvhetV1UA3eNXHT6l8QPEzSCFItJ+KAOZDf8QEvDFExNxkttWUjgOYLI3HLyjUQ
2Pvx1fHIlAKaleC8FRcmOxKvohvkTsWASjEL7UVaSU7rQnyJFJyRX+gDQGpqqQG0THNySxZamG/g
V0N1JaarnnicfreMYRUaJvqnu8Z1sSaURrH/+KZ4X4l3LBItCwhyinSAHkc5cTHG+1VMf2QsDu+U
qsDeEcTNuOGrTHSyFAFGKRf9+c/MDJldsyjDhkaA4YU3/vFNcCE3i0a6kUcxtWNFj0wENAcEIEAp
Ll3H8uYYmQSH8vncDPBXbigxxlSG9bsz35tzNfpGH7E8V5VWAJxKqyqJgTqqh1cHi8bfqC6jX8C8
jdViREO/Zfy+Mm8RAHZHZuLLzjhF5xr6bk3i5O8FR4n4nsIXgV0GnDo30YnVlfluWHhwCWjeEohd
OPU+x7ZbP9cO0Q08r1yudswG1PuGanspoU8rZZ/O67yw9rHV9xgSNI07HbeRFmgzWW95JzXN21kR
WwWLU/aIerdLdv8m86VlfcrMN7TWxq0LiheR4MoH+ejjCY2s2ujy9kas49BuwyYIUqO7hlxw4M1N
knDxoWv2PuN6of3fqjn6QWlEhnA2WeCCZP5rRkIoU1fOiJ49Ff/7rNt1NoXEIXgcz0Ne92NIL3tR
OEZvFmVdtPPwSJGP6KyJZtZdMwG1EBzwIWja+FTqiEtFtP8fjSP+yWCnL/rH0pWyFemvOX11k3yA
p03hMdgBBg1gRzZN1jpK5edOHYMKuszIkbI79seM3MvL7xwOEFZyErrnpVn/ijnw+qrtwB/jENy2
hEB9O4q+/7nCXzqn4F/++zsAx2jZT8RLizaOddM7GLgMP1RyDnIo/ojvfr1UE4Yl+YGUHJzcd2U/
u5NYFaXd/TZ6DQkbzkl+yP3AdS0ViO1qtmDC1cuWE9eRk/Sr9BZiLnaNlV52eH2M1RITjzqT0Tmv
Omb6Jm8vEDEdONNoUcfYGpR1Fs5VV/VakXMBfy0ZehZEYdmCIIUx//EkmUs1EQOianShffD8s2QK
GKqRTzcfDW1zpEyACWaeBpDyiJn2BECKhstPwph5dt1leHngPqGlmVPwQghhnlDaz3E3TF5NXAjk
h6OPnUY/rSfb+T/73LGUwn5GPnyG/lka5Meathb1XZ5qjofXuWrlAVNgT9cRdTcWdK8FnT4jRWsN
dR0zwmUmfx8eIfhFa4Bn6aIPQGHGhc4lg9RLWq4JCuYjzUPSt/1lvYZeWYDqrqkm0jGixpkt6VZi
R8Km/eZ+zT3CXM7dvwRbb7iz9Wbx8iPxXFKkmk/WxnBdbHeAbLvQxaAafcRStT25mLgwHjmw4uhh
mI6CHjp9ZHT/6akOTTIEFnmyR95XQjs22JERzXbQOaq7M2dcPEIWNKg80XF87hEyXYwFFcPPcP5i
nqP+lKep8zTi3sAI7HMnoT7dvSvI/sp0ZkxGrLCVf42IgeRNOrun7CZdeq+AoZdSsAJivsjaHlCq
FLwuTVDLO746vkQRx6QlW7gTJrIHa21yBrU2+j7z0r95WNRo3SG5S08K9Q+nXdI/VY5hDmCQYrCP
2eereZLgdiOCh2Dk5Q5KfdSCXn0OnuRkUIN0VyCQgToYM3EyMEeZwMd+upTNw9Ome8bqA6pUQxzX
h2y8/g1mgzj0rwk6pjPiVoH9YLQWyzELp8NNRLnmTiv2VugILzQygTA02B6+pBcJuiwkMZ4cOt82
96hHrTryqLbmdjxiX3ATF9alPJmyKpO7HykYcZIIg0xivCnaR6peySSKHnpBanxR0e8Vh5roopcO
2XW2Np+XmllFDmaaxdeVtKCO/JFBB74mkO6UXnk35o7lp4tP0+MlLO4rz4NV5NEjC1Yl7/3lgN9X
U1T41NBBUeuVymfP5jl3Ri8lbQAj9y2dz+Q3T+aIH3C1K9h/O26B2J0jY228EaXFhTCbdt8KUHnW
PMHUT6aLFw1vdUJDTooVPJ4M8EJ+Uke2QdNjzefCZpWWteC3sZqCakxul68JroB+AUPzw1+kzWx1
ejfhoMQsqeE1g2pd/J8ve3Tk9h4f0m6WjKEksc79zJH8KgxxWKnTUHVOn+XOKvtsaWahv0T+Tsmi
my1R6t/US0flldW726/2faVuWXUwWHrj/GwGqop+PnyRwLkkRu2hRAbOadnf+DHrfosBIu3lsvjc
nAPhUqKeEY6lP9TpLHjdGuers4QR+D763fNzmt8ILi7grZ83vq7qsvbgAKm0rhShmdqCzQx0dmy8
tmV8aiGRWpg6Xw3c5iKMIoZ0pbYpetLAUhGMp/Azq/mMuRmZxZ/ga0THn/sudQdXaE2BhHadtFoZ
RJ7Y8I9HrIurtli6uN19gWxGH3R4V91m1ptMyRfO+e0FxG5bs7KPBeWma5H+mo+xSAAG7/+HSEVC
hUJpki5onwZxACPJncAOUT3r/4H4vwuZ4bmePo+faMHjI4wzrw8ArDMlcvnVWcs9jnMOdyfq4tC7
FvhO/pkXHp6yGMvMlDGTGDkFxIM8j49lSOn30JG1cGk1F11kJxxcgbNz7zd9VXl/tYaWv1FxbGHQ
CQA/lOu3NYRG2NlXYTdj3Xw7w3T+rtuIKC5ar3DGnUEGjXdx1KeGsLUsEA9G5d0ZeJiY3O9w4GMS
LUDnsZaifX818FHrpc1RnKHnTtdb1ynky/iHg3nNnZh5uUL5xrYzMKvTM5P5NcwbHLt85FodyBht
tEfF/1MgZmpw0SYC6sErelsxIi2VYDb1hEhezYmoeD+FSFXCDPWCPZjozfOhWtG48uTjBtXHBfFx
vGqMOPSyJWnNeNJjCH1kEP7wLFITSIqd2XdvtjNCBlfEeQIxGYZeyPQ9HpogFYaMRSaAUL8wOl55
DZ1MCxHldiZH5STjKwuV3Frq117HYb3xWg0WbJU44JixxsdJGqmPofnWftWLX8jdZ8SyRomI7nQb
q23gWfONTewUhFbkcZtJ1T3kYlaxpuSlaYc7JxPHok94ZD0s5GLY0EmNnv1mz2NwSSvsyaP3Fegm
OtOTguHrVIU6Gi8+mSeFvubDhzWuo6M9aG94edxTi+vFx9obtnABhu27Nx0nmPm6csvb9IcrIHZU
3z9nszHoelvCjAJs3eYUvrajT07x+SJSNS/R7+tsX2OX4NCaYYFiSUEehhaoi48hynHQhcLqB3UL
JWcmLTMGRxM0GN6XrSMdeRnwbbZ3z0QTu+oe1CByh4lIrvZH9hIzImhB6oJeJpbfmNsW6fOMsFd8
2VKS5qTsVbhfalUD3CfgWSsOfLXoQhAu3VOvs3x0qW8nM1D+Cy3rvLXmfsgCPAG2ZF5A545ADxQ2
Qc/vf7EGN+pFyCgLQtaLjkJ4xXAgmifcQgFag7XmInB2MBuzqcn2MYwNqcjxW/fqGMUFiEIp5tvK
S5dmEmB3ry8q/YZFNJuhLKSa1zw4IXH4ZW3GuC8k2zBifNa4YdLnW5IMx2gLsFxyd+azwyytUEPI
ZEqsEtUNUr9V9rD2v55f0r2bbyLgpcZsIbPx0i3Vf0bQjHTLiShFbkidHoyDrat0vxH9U3jUf4JW
Ki+dl9s+TI0mXH3M7AKMCOdY/1xbHYV60pN8QX4NhEWdIU+jSghNLQ7reDEr0jFlM+mcYUS9S0qf
pyXEaGmKQ2IpNxG7n4MmCoQxmSiQQd8l5ixldGpJK4GYHvhvADFCZuEWq6W+6Fok6o9CPBXUNPG5
j76nED6F3y6cO6krUdqIx2pf2auoT3q4pkCfDDC1xE51GQPlJR5V6/kB7WRgzJEL4sqbXxXCRd65
XkmbmL8rLeEO76P0TZ3VAwYCNZFnQFbPK06tNh51N6HN81aEuCPpwsPytMKAq5FY5dq3G5bjgcTD
LqM36CIVC2Y5cYLwVDuS44FSFsA1Vh7wR/iMLOUWcICRoc0i9Otx+KG13SSkKBo7IpjcBcYPVCRR
PjrhGiv/eU2UxecAzpcYw/YVRPvua7kc0scP7u6Cxx8Omeeou6cnCoqgPg8l04SBmnRKXgaTTIyi
LDxUucM4GtMc3r8MOYfm+WnABb1Z+6D1J8k2z5K927j/Icj3Vf6igbbPD0JkdD3qLaLaXb3eKLQ1
LsqcvaZNoDR4ZHfMCoQcEDEnpzsFXPuDJBirVfDFpjeSwJrX3KXdw6kUWhmVxv6inilmgozeGwCn
Ki5K7Hcz1xjYv7/ZFF7LM4MlaLKOZ9957UfmzoPyeahXnKRhjD/z1Dwyk4fuA7ki26B5VupRIlGo
tbBDLdDLfnzUXtblEB9isybNSX4Fgy+TsnklXuK9oLHcNPYSZ2cLcs2+LPytNRtHGGgajAyeq92E
fN70QoBJS8dR9GbgtjivfZ4MKidcm0nlVWpQlBu1lRlmc2J4b9FrEk2K88ZJAE33dYLmejIFaDUV
2H8ubQNYx/kQ6JC9B/GfH60uKbNf27Lw7nXcqlXtH372Z/kZgn3eBI5O6rE8DMV1l59JmqTxi3IS
YWIklU3cQcFBXjDjUoZv+eTtNui7rj0Scyb15rXTMTPZpxtWhrqqRGl3DSfg3hdZ7NyyCmNp8R/7
xcrHS46YfT+GZNsaDowlAAfm73oVgkTlC3V5t4/yEsKnPR/3WkaSRfQlTio4dncYNcZ0DARy60B7
MGRmId85KLXiHlmTvl6v911W4Zyc8H+eaYR7wyjqlrY2ejg7Dof78TRbM2MoijAdP1XcqDwGbxAt
nycEJvw286JNIl2Uy4xgxv81Rel+sTeBPJIqHnpz7ukrbYTzAdAaC5GfR7xhLyq4iqvBoRHYaghV
ZWQLkZJb25gbXeQhWgA8MzJB7Gd3e73NCLMsrNfox7lnk5j4eZTtk28rxAlJw7x+Zond4DOyenqK
V7arUQ6Ctz4nEoPfw30NWATfPtBKY78d+nSo/vEbD3g8PQDpQGFW4y09tEUIprbIMhKpEQCS/F4h
qmB5N4FieXC8Yr8gQfSd7BW5RUypjVu+qQCjEL1vJASaNIncnnR64gPxQXdFivj/EIBmZdZWrLA7
iv+BOZjDRXiAi4TsAs0ZoeclMqGwF0hInxY/Iw1K3Y/0evkj0ucHs8P64TRZPlg+vZFGcL3yyPM8
rbs8SiqEz4k+HV2vaHtHdl8kx55+3pAbr/pv6d6iy4/OLDM3rUnsqcGrK52aC9Gi8NY/sNB6JYtq
xpnXwxbhSF2MWDGi7iXzF8gWrwpQlH43IWomeXe8jAVYBzoeqKBmJgbumV664YRmHnI7weJHaXVS
yoReB5YG9xJhghKcY2nAyqp1BQTAPLhHL+w7d/i91uItyENL+CQt3gYu9gQ+hOIGkuGxWOkJFMnL
fXHS7DW/Ypb9nxgtRlFqQOW+ikX7NaWDdWTba/r95NTuWACI63xPh8XUtt94f0x++TZfldA/l1Jc
vQu/yW/X0nzvheOifi0GqPXZGdtwU7aXcFC40KyoI5EgtieXWb8lGMxq2vjFBaGVijefcZe8wi5a
UHP6tu7gPQJI7z/w4Q2sivLvyMHwOMje9ROmAnr0sjUHVwyWlawaQ424TH7jUBc9hu1alHhHDDcS
2Pypw8TOmVPLG/pxvfm+QrAOgwPDTql8nHbPYv8w8YJ6QMR8CgIucgbfH4Ic5+3L40twaT3NwtTw
YRzWYDmzFB4UI6j4YsOrOaVlb8a3vuHBHp7SOqlcq1aoakB8vAdcEpjPG8VjORyMCwHcw55WTW91
gMASBHC58ZsqugxtJs/KxywGIspA5PC+L8A47iGaJDaIWk66jZk6Oy1HGyJW8GfYh8dD7bf5QsOS
Mgh3Tvra6rFyxLfCLE/Svyv+vaHW4Az9KFa6992P+zOnPwX/lhAV8XsxqpTBqDf8JvdyNmQOAOdh
1i2n56f4Z1ByFMct+bJxgqI1tkwBCD73POZqFzj9LpYNiaCw/VcNxrD2z0FMvZNzV+SUjqqYfAzJ
11V6zntL3peVi1MpxlLzrla1Cz0F7srvb6fFIY881MH8hZApoWRZB4R3oyAut/aOAQdi2Dwl6jIQ
eeNIJDrusVjfh8xpkwls4Ud7wdi6yrL7QBeEk+2bKzQVUglt0DbVJpc8nscH5/5vGzHvujdp2JDw
2WFvcHflHwG4F+LujmoxDppow8BTLgvjUrhqvvGDzkC/hRcqxSwOS//AJ4rJY5O2fuvoKQu6mYs8
L4+WlOUf65AYNEwYn0S8ljlb3J09GNI9M/WvBVXYan07VyDvvxGGoyA6Y4H1lFRPg6p8o+nmGukZ
lPjpkNyFtnvKT7KUeIo7XgDBw7nVsCMFMJiya5HMtFkI45j4fmk+OiFJbo1/3/GScA/ZcJp1ExjO
4Sk36+ZmS7V8QZ23S7XsVZZWmLWRprZRTm2ZH9WsIgLPw/EH+Y9TvYJsomMwMymabdditOnycZys
UNoOTTGcSbhagN56eu7pu/TWOErdQVkV1c9roz+Td5GDTw5Xx5GOrMsvxfmMT/hghK2H/rM7fqBF
rVhbbS6X5Uk7wsCAQXsr8LQ44k8WTMflBpjEIfc+ewFCfzp7lkI+cYWIoxo/K4YddQZnkjkIetES
YgDtz3uEBJ5z0REY9Np6l194uvuGwWH/UT4V/OYsuWYLNUnukZoXEjHBoXPwswkZweGzUc1ovFBt
1z40OS396B2mxeODGkFM2IpesDmaDD5ERRdTmW7BqTgSsa43RY4ImQTOlaLv4nTMDxjbaAVepj2C
xHFJErFhd2WTDjhn4X3odPO2Kcv9yaJMkZiOps0pXIksfQsUc+il90aPGqsbWnYxa4j9yT4Y2eKS
KJVEtokhA+FJMMUUVO5NC0R57KDKCTsurJ9sHe+8jbbOvAcTbmVsBGvyFS9ronPTtnEAHjW2S7IL
CQWWDtTx0PXcqW8pZmearaJnyeNnNoOzi/6rJuEfKJEs0j+AU9kNkeLtcOT3Sr8+b36NzDjKcRmG
8CybysXvlDJvEI/xcoWgCM2aNN8SDavYsbH9TcIpACjWD0necWhfnITipG/GZuRtRrZff+r7H5uv
Ks9ZKt9WYNWNNdT3jrzmI62X0mZq2V1Ed+s3KCpvBC/sVC0IC7oIQtFUEcPu3CmZ7cbKFIPYh9ej
jpASqqIHND6wr04gZUecTeCOE001pZrVaM2NAujY+9aJnamT6tMU7Z7mJOZ6diWqZ63UCHHyWwss
S+EJwIXT9YvpMDZKV/byS4UTK2cA2dMlhFFDRpQMabDfJ1jUtDbPoxYX/EUBWZO6rbxaZIG6KC6Q
IFdonPMU7tFF5yFFeWOgI4kVLYi2Kfo/XeL7GfNXmnLlEvE49tfaoh7toafmnmCbkbVFZpGcJbYa
/z+8Dd+J506CjnQtUQQTz4/maLx4P9dyult7rUTkmsKGhAJ/EAKN2DC0k6WVFI+fSIZA837Ry7Up
NWJggJ8lRKn0R5BgCJKfTUqsL4D+5fFVWdMKKMXot3U/BbozmIi2QQf1neDQol6kVSlSm3EMMMBn
JzbFXpb1RQVw7ym1dRHIYbqAchxlkxU7uK1nlZKhDq5i5sqWlKdw6A0yTJgU1JBtENbjX0RgI9z2
2FgpzktIRvFdByQGZPgcp/ySwkdCtUakDtECSSyuoF5rgsUgLjwEGi8NtPelwrQ1gXR3E7vyrWSL
F9O/px+kvErYGEhfih/xBQ5PcahJa0V6iV5eQ3EbV9J788iqvDJKCIJ4VusZo00k3OY6Oswtn+Cr
pe+JPqQCn57963oZCR+IHOxujmVnm/i0uNeWtJUUsd0SPZy5tIPjtHAqbWbcInnRcSc0sADHitAW
drI7VAwwLYOHhRbrPfoc/QL0RCcFzHt+aDme7jEWJfMLMARCagXxxYN6+fPia3tcFkPO6JX3d5Q6
twk18OIwiHRgatE5Iwh7MW1RlT0KzFQLX/8etHeVFuctB29XE7SMi9HuMNs1smNTW33CX4UxHewQ
+NYBiG7WeaMN/7ZYuAFqbBnXCPQuaaw2IGgb5YXD6feqGLMDi8EmnNNIsbE4udUCqBpEv62MXfZC
cLpYKcEIfbnu/UqD91Gtm4H5QR//gj+AMmcHEXkxTldGK6650U4GGl9tdukxG7NyZqh6BnEoZaLJ
HXU2DD1kKsb6q9aoIHf88TZTRLGB70NOtw7oXCoCfT3gcr6zFG6SkapWVRDi/fVgglJbEvJhAQoc
fdHZBQxr6b1QITF+s7Abz0V3QK6GSNGETwPj89+5AbJaHAPxjT7i10DPXXnPs+6E+hGuoe88OMHk
KGRGK031kpq4TS1dB2Fsvpk4evsGNKvC8hm8FhivytHBwGPK3k8i9E95/nhqEGCNGnJg6iT4HYak
7Z6WSIvO3+ijJMSNLtuN1x8EHqoaL42fFBCNw3gpiOkD1GzyitlIg0U/REo+nayxG2cMEgT6533j
KCbaXVOG91anUZDKN33e3i2ibI2A+jPjfzEBLVmajhl2q1p3WRAisV7XiQ3wZsZ+1tliZqZIL/p0
cm1MsUYpHdCIWcLJ1LQo4P4bw1Agiw619C7zRkhs3V4V4iqXtRLvYzx/d5wDftK0JQ0VEZqCzdjW
c3HzJm+nRcbefGWJ5lJ6s3uaFinDixJgWEDK0mIx4L4zoud+8oLzMUy87NsER2s1doExRM2Um54g
Mv14H14bNNC7voi8vptoX28Yv8NSPP9g5fs2eFey2Zebp3dSayyTv54vkex++Am9kX3oSOXPtzpb
BhNlv6Ki35RXKF8/IIo4ynpiomVmLSAv/F/clhi+fi7yVFzP6PU1YxL55ZleM5o3IbMMlBzKCa8t
WSkM1F4t16y/or15/cEs2sXAJLXOYbINumubJMQW1x1MPcGxUxT3n0KM4F7X/RFCU2CQGGzwXB8n
Gk9A2MWIM9VXbxApOXGlVLZiW5OcM9xR8xmJ8hsFtC1vStWdJzlXQlzAyKaCFhLTEY59MYcrGh3c
5kx2+pQnMmjASHbF8U+XVJiLwJfMqsc77X42cuK9jbAccoJZV0pFRZopmlSGRPOtDgEcLwrmZw2i
K4MP68/HGEYOSNM4ePdRKBj/f5ZbINUAnWYjou2PHyK+odfDPVyUG2I9XlHYeXRwyfqoIDQrqeTA
cKEVy0rBTIwDf1RBPJ53jfyuPyqIrq596FOWWpYIfzc4TGP9qxK8snonEKGJavcSfgFuCCzNrGZM
0zwI07zomC0af3PkcsI3FmtUJtcDFY1sWZ57SfuWoeqaE3kXq/BJYZTXFK/wRRn7YIN0KCVUNuO5
wFIuVQTAzz1oopMwiF84FyYz95M50kM9osTQvfsNiTy/88g/jRey5k8FlGiRWKI3QVB/79n7f61V
Z3sh56Xir4ytHSHzx29bA6kPpPZNlEdaLSGthREJDBsNcIuxjXAmAMxY1rt17WNyBQVfMsS3Z3jz
fulM/LTO8zclaIDO/zjoV5pJcf33CPFpP0Jf1ayepqRkGGXkTc0KfiVuwnpDCGHvk5pmbv3ZGroN
rijiXxlCN5nXJYI/+KoxyU3UbXK3e9rROfwlmWO9WV35UH5IyHX4IvfMGSvD6gJIQinWUTdBorXp
c+HpAM3KQOPbtWtiPVsyp4LKkmX72x4JYClHqq8aENkAnDtTkGYFPsJj75QQUFvTlo7t5brp85uC
BU6WfEOar0/aJPPmO3TZkR/7htg8iUA3Jlg0hPdtU5SetitX7WjQR4cD5FCAXoNQHyhQ/FG+6hix
iE8kEHETlXlPSWoc7/1rwGVkfLzjwPbhcBLG4aUHIISo5JvBMP2War/kUhaDz5n9dkb4lNLPPZl/
UJX5tAv8vAYHUQiTmnpll6tAaGBT+VxoYdcgfWnz6MdCINdvHJi199gnAoqLA4IceZQnX/NQcC8T
LnmYXHDKGJEVXnkh08RdTprTOpx21BT9ic7lrIGcAin3B7X6lqMXDBxsIUrX9x7J8HeffvG612vW
IslN5SKqzD/11MprQQ0B/tVRZBCnIKNeMeZWW5SHZqR67Jax8nNfPYuwb/8kvCwC0X7FVx3Dev/9
vCy5f2ByvJKwKpAW2nSp25mwwshXpCWNmKlyaWlWK4SUzUdKS8Z+ZYoiR5t7WGL/bM0CFM9SqXfv
ZgOsc0E6ig4A0gLB0nH4XeggLJr6nEnms0IBe6EaNrqMweLsfoHoO/2CxND2aLiSgq9oChiu5OLo
gIphV66RgMnoupMVC7jpfuYxdX3xU+BahH8xO3DvADXTQS7u4Bld6ox6LCczR4oisDs/M5BdOd2M
SKU0rm7E7F9saJgKrxXh/UXFUFtL/PCPmVNQgavrNURHugY3B/aa/RnTBpjh3KlKr+6UrDTetWeu
2YoY2ZJtGFHxd4Qsdfua8dU1eCWiNue3wT6R61n1HoXGdHyForD0Z3x7NGUCURBTjy34Gflz5aSn
H6MpWWFs1H88zfAJ9iS8b9Wt/cqT+ffAFTfE0bfapTN+u1grOrV3tk2UFjKD4PPDqZ42qRMqO0Ac
yPfwy8TBEAC4ejcL1+r7SAPzG1K4smI822Yt5Z8tJGE+eW0IGDyR76yddz01LqEcJHrgi304pMX/
35Ughnyl7cm50On8VcPz7WP/w0c4L9qUbNRDNUrz6SRbC2nUn/BsXGl5P/sSy9ljIC3+wJUk83Xn
XdrrwfqMg1ZB7Qd6M39TTxB/B68AyBsLWZMjOdmwt83w6+/5dapc3KfHUD9z7SxG7HkVHQF2i9cY
JQxEDYwTLAMBFGAwRbWN6Y8nF52FSfMEOn+7FAYSh6HLbF7U1yn6xw2D0yD5zdrX+ONXltFyR23R
sK48wFy4ViZAzU7ynKY1HIqtc8+6+wyNGXwHbK+AW32spXsbm4AkSwjN29gmUFsQg+LfMx3Ey5+T
2bBo7p1VTWUfR3NeiYGgTveMAU/UcxDomm/noJAh9C8lud5nkoui6MggFx/0VTMzvKhhpodDIfRB
/hd2Ym/ceOYjKiu1A/slcx8Xnzu6sqYTSZKscrSaMxeuKP7kySruFQ0Txeya7zvxhox+E6lE6Bo+
djs2F3iePFOc/iQ0Ja54fWdMBRrvgpRO0nCa5BsOlAV+59U/6RAHucGPZ3xBS6ugH348+y3gwsEg
C/mngW6NZYRefEhBY+rMjtEB7tzx+VKZQzVJWx9MNvll55JN7hVyYCU8/nrsvgGRIqkZKiE0oBn3
IL+F5H7FR0IVfB5bc9p16RSHzp02sA1jlfEGdqLBeC7nmBv47kmHaPkie+uufoGIeugY38TN7bqQ
TG5qjbx/OqoKH4QfFOOKRVFsIyxhU1j2HF7glm2tMyETeOr1dz2iz9c4uHlUrs1gfntc6DQIrzCj
0jV5LgNux5cDC5GrNIhLWCCPEmrRjEC7bN+KLyYgVAOXmzWFndCWx6E3zGIsBztWZwb80Kj4Gqwk
4zSuR0hBq3ADP2xZYTTqf+sBrxVoXeFjNY60YJv0iQcmtZ53v84fM1wCojK8N6L2TTrL3/WRYEf3
rpm1UCU9p45TlTrrt1Z/dJUAzUu6Ts24Sg/qiiNodmIndMkiXkBLib/yiu52AVGg+O2Gulx1G3Cw
uU9T8skqZCml0j3J/yiVz4kEZgOORq5HBGa35Qkck8OXC0CLds9M//Uo0EKu9eaFj8TD4U7chiJW
Ft/RSxIFD/o/0711ALW2v59Hvh+itID1UxUmWM05YQnMePKG9SlpnzgtOcFzUFWRRQziI6Lts6nf
do4u144M7uXhncj6T422D84XjZQ31QIpSpbw4w+EJfB6nftpIKiH13wfegq3VxdYhJtpUAqUeEUy
Cmzq6ch/nECYtIyhCOTL/gqYRgz5sqdFN/W/zuqJeV9v4nc7Qf0dp4hpi5bHPkDV1NNGmCU01KlN
NVIhI+b7aXhA7RnaVPCKaUStci4QmtvtsStVc4C2IcylwFg7mDeO/3tp7rgrKebpUQ6f+qRzifIk
x1kWGnMT95T68X9PDJzTiEmgBVIlEQskJ//4dd+pnW0NM9WVUvBXmOJSJ+bbUi/Mx34uid8418BS
SQ4eYQS6YjqGudoSQhYRmcnhGDTovhEx4xsgZvx47zLUqpDcvC0C8DJ5/OR+kRPCg24pOgt/fOWI
D7TQEwtAEB9sVwnygbHN7Uqod02ufVEB+AFTnhsJ18noa9lqGQ3y48KPNdTkG/fiy1yDDvV3IDVt
3SPWmtLcZfw4RHN6TCzzGEIhrQd9P+kfco6y9D5AXIMd/xdVJYxeSfqHN50MKS1LHdWDiKuQsHDX
ipIFLj5ehS4P1OwYrio10MWFgOr6dbCK2E+t3t/Hl87gd0Tf1K7CfZLEs/LC32x9QaRkvR4flMVG
RO2yc4JAdGniehJ6SmVdChO01XPv3iLPH5SWKxV+yg9OWTHkoOUpzB+OEbZ6CPGnHFsonhjnsYRJ
17/yY5onJWFSRTZhlv8X38QbRGgU5l3U4ClNY+HTFN+sjqhz9hm5M3MkJJvoLGZqxaQvao17UVTf
nP44xJqqSxMx45ISurg0hXEa8NBaePOu8mKONFXpcKNjpl9Ou7uYSHSGhd9ZdzPCCakH7mvv0wiR
0pE7oy3ElYV4kjziJq9qJiJ12fV73mbUDu99DEIiQgE2v/UeT9heeg1aVUsWuDq04uA9E+jMzWLk
gUMNe7+ysQWVc3qDJxfmc7BP7vEzgWf9dwYEyVUoh59n06nOJTUulYzMVOrv/+tc1zL1/+1ymfJn
rElZuP2QGuRG3c9QwnUTOVY7DD897fqIW+cXJnBuCQ0WHNatysvP0j3n0o8+oDbN3rDVSoM3UkOr
yLoBh3zMyWjymN/cTLJRrYPeRsjAJ9d0PJuAO+5ngxfwk2DoMSaucmmIHD5zTEjojvIaBMgRoruR
KIk0XEPpDqvoLUMWKpXADnjHCyaMpcgc8wa6rqFr6/pdP9GfedOZ+iQBUeuY/wns5ipt70OoClxE
Nb3BDKCEB3A3lUWmWjzpnSNMBzhzoNtlLxAaP78UY9JaSOGUOB4Nwmrhkkjq3c9ORQ3CL6xWMc9c
Yup6w5uZTJ45i3m76OL2P6ycw3Q0ga8GIts5N8XQoQcFIbnMRbwC0aFJdINuaWAaQe56xop6DPXt
0HlhAE3Lolgy6oyhA3Sy7V6wmCKG+j4w4GMGcwejBgGlT/7QWgrQRBmQ8PW7GMvxNsUmvyMZig7P
tK5on1SgHoWY5CoWA9WpGZOcG1llOyVGSt4qewkpUyUGW5+uQiOa1jYNWHoJN+LAsyj4ylo9hnZa
b6r7QDErv/FXzKp9DvfuJoaqoGoPjmh6xSvuS5BOoeLCxPlSGHS3AC+AMeD0ai6ZK6nxyHKW2bSV
95jSfgBS4HMqlBm/LPY3nVwSEc9LcigYJ2AASt3cUjE6IgYDtHjrFTGdxM85m0f3kCY2Dxrvr0CG
8nBnEh7rQGJRQyMs1K+i6eYvLOmrwcsJMBI/BVHgFXb0wh9I4hwVYyjUFa3Kju0RGrDxbgp6tcMP
114L6aS2vqIeiZ4wmk7hKOnzDd+hIh+rRapl+EDQ/r1fCG8BGiDjgEwbuwx2CCzVEf6s52oeziia
j8fnerYd3lqUYGbFGaEgjcOwMHAoSGPjByRohhzsnIMsSmypdOnOtB70RtcmF2PrM/nszGqPMWiX
7UB5VKlFuGtCiKou4Imh/2kyu1v+tJ9VhOMbbzlXV39f2+QH2rMSabheg8L+DesGxtS3eNDk32th
0fPEG/v8pZhcDWbhz8NjUJd43uYUEMcfsNHKpR7ytU+9yH1tq7Uh6ReU+KpB6OIXYycYyItXxP1+
8KfkhuI8/Jq/y0XcIhZGbr6gQIZJfZb9bIFml37oBc8n4aZRHxRGlpfaF1VTUAJCArkAu47S588Z
R0NI+KEeN5/yAu/0ItfTvxWAhYg5KKwddki6srPUl/BJ04EtAierF5WVTzEr5EehHvzX4N2LLgDd
ugvpAb6Sxk83/5tMkhOdv+W4Jjdwros8egOcOxPhQGW/4tSkPxsGetv+XlbX5DTLKHicNpWtqF0T
P2R7KYgK7uWXvVPYy7D2069S+liI5DjVXHHRGMSNbseoIFtoG2nQeMoDtlNXVYYdbKUn44k/2tRv
DmVzhPHr9ltEZ6+Da9cuCyuDMwX0qDtLvmVNd7P0055A0TKt/QSg4AolQ74Bp5UP5YJ+38hfzenO
9wOBNR31GjL/wfZRtHTZsKOEo2u8bxiEP1Uss0Q0COGY581c3Vl6pUgl6N+wwk3IvRmMR4TCzVUG
q1ybxMTwX9aZDZuoMRqsNgn8kGvDGU4Z7jVJiFTLYW/EnaVk8VWYEUphE5z/YPHzZdHDQPng4g8F
0ZDjB0RGktDHMf9CABazM73U/JEcHxLxNO1YWFqbKmTEIndp30G1vP0GAEmXHU0KZXDLYqxJ9kbj
/Ye0HIs2vjl7kZFvfvaxvJWYr4+O5hmuvfq2I0vnCHv8+VYmjBudyNeG9Ee0slOLWZjhigDLXqHU
5ujSp4slQS3UjlsLzAb6SzyYn/eeK3Eatnw+GTEty5X7fDy5RQ+/AVVS3TsqRMq/Ki7YWhaSFdO6
32/3dzK8y+0Ylsnst4k+211LGs7jeTT1js8XdE6Aqj97/y87+utIaOV/vV/lOmbfjM5zCYqN2HHd
Mma61UCaNw6s+fz8VE+TekqnjyCiIg3I5OtTLRAVsKpm/iPitBTFYjmoHfvi9ubbexwggDAs6R3n
GvWb82qe7goQUYmYeOZYk3uFH13CFWy23wwWZTE9ko3SRt2hxjGh8p3/tBRX+Dnf3PFQuiaxfzGt
iNhX+rlLfZKLAAvrOsCtLisFzzSqr58V2Ae5ozjMKvfWNQR95BQQx++mu92gkQH507cajtPBwV3p
AU3wZPF2YgvQQV29cKRjTnL5tMKpV6EGncbaw8TR2s662xO1P2jIj573p80hpfl1rmfPBui5POwx
UoCOn6HZL0Kw+3wM5Yo2X3L3sPmG7PpqocASy+OMdCeGDZL6KtgreyClIWhnmun5aNwwArh3Z7dP
Jlm/vPqcUHm85M9w5p83WrTo+FYmWLkxQvNZWK6agvUuj9vFtYmaB86Ll4gohoRgaYYFbgpyXbUK
CyAVe7uHZ2S5zG2gV37YimDHX8uRnjdjLud2sKp+4wUcHdvH8tg6BnUAM5YzNqpY8J46xubb+LKb
0mbB/vecD6DA4rVqDCJuu9BYeGefum+7KqeiOVWNUQ3ysbqrxK7UMDOhE1hw1lMKyYWxMqMxRyk3
ltOqjBAMpFqW3Eb0gxxRRamYALTH8QmenaZtRKeExLfM+2ypJCxCK5hJbyw/qeA5rjAxL7450pey
uIyMZoqtYw+6XY491oI6ksNjy2OhjBhRvsN4L+vMsJnP4KONQuQO6msUMfWTTaJFR/mH8H/3Vz30
8/hy5qJcGlpNrWI1R18s0HsDtKBN2eV4r4wyjrgqLNQy8i7LP4K+ZJKJdiLmuyzFgRIWBAfHOdV9
eoXOZ0rRqP1UggpZfH1I2PzQNW7wbS1qgQRk4U1bjeRGs4ypYPidOSiTWSN6uXVAd8NYBuRamqh/
lO5WNUOKRWaPSS8W8bTe+0Z5gv66+BcsYy0+GKE2sGrOz2pnQK8p7Mqyel9IhBkraS6kcsLSgqCb
fj68SnHcbi3a2fFQuwIKabduzYd/ZeFMgtUBqCaTyZLnAV8L29Nxj+0By1igMT43Gz7lJmQ9kJ1Z
n0IJfZdpc9/MVlrDhltsa2q9pWeKHGaEOneyg1EHMF9GNkZ/6ka2+Jq/ohlXZnjPDZoLxIPdCpB+
2unYm7YVe1HLB+9fM4lvV5SVx2vijaY5kMkGbi0GEa3H4/cd6QdkGIdlP/bysSDSn32rtFo55sCt
/7kwAQTCfBk31t8lf1dhVIDB9YFbwlOqCjvvP27tIYROLpaazzLLsTQwIjZUztMJ77zXDk/J17/w
nuUMktUAxE+1ycYVGZRJh3S86i7nH6XHuBpGTBj+PG4AS4DnbniZ8xYRfFA52E9YWHc75zYOC2TT
9+vxU4Sobi1GagVUZsTVXV6ISrt0D+gfWwmyMqtP6Ze0D0+iTswuQdPNpw23c/rJoiH2DrjNVyt6
NNERR0qpqYlcaBKYURvoOeXvmySpO9I3/jOdfMzDNf75BN2wJcJr+N3QzCeF+9p7/Y1GuNv/ldA3
d1joTfa8e9IwhT66PUv0pGA0sKOB6SRyj2lsfO04u7EjbLfT/AX2I6FeC0dllkDYKBFylZWKSO5y
k2IWeMKry9Sg1JKDNFqW9IiQSnXZ4HF/0b3WRlvMCGVGRoy8SsC3VXco/LfFYUTcFj1RBKS3MliN
5GDyKFNwrkv9jWgCHaHQA8R244jVI4X0IFPb1+Gl/+UZn4QWGjXkc8025bsqJZ9BBYu0p/vulz9a
pUcqT8vzc+5GVxEasamrPiY8MnLg+pjixvT6oT5hCYwj9hNibqCwbPjEIB4NFWBj9qaFAU9T3/LH
9h8fEq1BtpQW/oYfB0Tuunl4aFpKNdwL+tvnsDh4gtMhhs2Pg53EMZstMxZU6pm7zkIbQth1UfPE
/AKpGOUflUi8zAYwwgKKjntAazbxILsXHntWyv8ojEZueyFNVYJW9Nd7OdKuhFs3zmElVC8VMT+y
0p3K344jsdcX8t99X57ilibUx4+jjNidk4iIYagm1hyMuOGwE/DcCoAuJlODy1UUr0E7AZ/KuXB8
AIi3umnIGEqVbtChLBT3l0Q0ac/gi5iRxgJWEHzKloXCEIKiUJZqtoraMiqTHc+KjnzM0mzIPNHh
66H76nSG3R4ap9O2gTXggfSDQTLm20ocg/q9Qifx2syLX/j6VSO4gnnxIEa/djDffGofoeeoggzK
oZ11VpmDsmodoaWTTLYWQavklvMm2dw81wD3D8OazhKjBbCq7tCtMbmIQ5hrYcQvkiQUarfeUR1N
3pehbS/7HH2xEIqh4xtdS+e4ctJ+DfWkHgmQUg7rkb2vK3Lpw3WLsgXWuf9Vovq06tkcinXT+EKe
2cVbV6/VPfKmDRdogctvN7IIFc5PZ7wvvICGs9QE7Os22AcIspwQsOZEoPeu+uoKQCL5LCj4NEPh
jfN+Pe6qtdH8+eHyhfaCapp3e7HcWfF4PJDQTjng3iGJ/nWpO2jTlDDRe71FFkqUcXZcnEk4KfTW
TRnhju9EokRoxX/n+IQq9u7za4knaOr9di+d4iprUXFlng1InkJ05lUtBADNqyXnIV//8LU6wfBS
LKax6QHXR5p4e9LJ78HNwWBsbU5oAzCZ3lPBGpXGbRuRfj3jz92aNJiYF612/YJTmtTzxach4v+V
GBigKDEynKgxMjdW+JMsc+9TIftVUxHA+znFZr5TdLYcg96TjrSahiPanHrwTnULo50PV2GsqlBZ
/yS+lmjaO3ZUj2lfiYgRWaBPi2YeDW+KRqcZnJpTzHvBioRdO7SP/vHaWDO0nqBCWwgnHhYg5j8g
nLx6kFLMen0gxglwo8QAG3CyS9twV12FwQFIIZEpm/1iN6lWVk35gwmGK6gGnWkWznEXkRctQ8iZ
H79FK9Pb208KVfbTNeu3O9owJ+fJWENk0HIH/l3D5uIw9pLtXBCW0951RMjbLZmaOQx3WLUJ1Bf4
GcyyOBvqRalAIVQxxaxufkKEil4N+p6faXVqOgwhhEbLUx8bos8gk8M42o4wRNRx1IfS949FyiLz
w22XvhDyOlaAqJewm38Nn8AVVGQm7Thqk7LNbH+G8ushMKHH07vGD/j0tvkQL+potHmVHzQsBJYD
Xz2f7na9jncnREGFkw4qEjvtEAkcgtqvSDpGsCKfB81V57yjFilQWjvgZlokHJqehnIYgD5+OsjZ
imcjc7vpihdFK4n7psxEz5Y+fzpt9E/cy3Cj7d7hyzoAcxJadWbuutttnzB/GD1DQuVEMf++hKJX
4Vi7ytJJdf8itOKOmUAJaekCHOlsJjhtje3O7Z+gtnzS9Xj8/OLn+Ts9ZphKs8kOmZ3poeiYvJTE
/um7sC5kbkBtOr9pVzScEoqtEx2EuSsmljJY4oS3gx4DYKEhr8REFxkDp3C4wyOspndKGhLOLMU8
EIN40+EXJ7ToS4gDzoFjN5FF/Q5cKqXVS1YNRkFiLHtVu49M1s8vQHzmRvW1NrEBkbJ2FkABXW09
HKv7yZJ5OD6HGcqP3rBw+sys3D031uRoFqAAlhCnRXUu65H8AoGD2OUun1FPhN3BurVMVQnosV4A
aWKPzTvKj3Y4IaOuphKDgEhGiQhoG8wuP3FmhofEmV+lQ+Bkq1GvbCRtIyUOdCUNpkuFbNr6gqRe
dCQiCFeuV6rdAlUdyS+9R/DpFHqm5PUDV9DTd3KFejmgEhbgBjUxvzY1nu4+jksCWtacVLZ57Zfg
aKEBQX53g73eFWgBhKAaZlt1Yt3XPTb1ls+ITPAFSpGu/d/GqXhPons0CnuB0UwU6iGx+y6juQ8Z
aEkfAQfUU3L1Si9ug+5Lmi2xrdlxSdoIhe4+WmEYLeyXWRAY2Ilrpeu+JoWnXZoIk7R5/M+D1AZS
ytxF4g8JMBg6ilmb1+PZTHiwCiuMWd6b+AQB0VhOf1rC8p4QZCiV/Zzaz0obzqLwMM+V6vzyCptI
rFx/Rnct0Ow0bHfD7zOqchID+GFU7GmjBIo1RK+iX9gPjOZwE7oxRxJEvLWAjByDZRtVwYzmSihS
AHFWoJ7BqKfmALhzhJZnYq7cNM7inbCrwtdbIMxNPbkva/xO/VYRFVNA6ddZ71eHKWTlnIoCfaPW
YXtd1fpdxeh5ik16BcQ687XBUATHiT7NsdahkA3Db9DnJ6/fW1GSQb121TLljELZ/VWn4WMh9NzQ
8KbjuFTZu2n5qPJom72zYt51l2lvefYCBZhmuUEKb1KfW0qW6AXEUZVu9Q+NaOQu+N2pfWQTFsNn
MH3CnpA0KjRSCwFAr7RMksK0xbWamJw8rCe0gfyWvfUJKglVkM2HnhiRo9y/ye+BpFOfSD0BXVml
Oo29HkJR9HbDT8kUkiLDkQveRITaEiG/pYtXAl4aMnZrMd0NBQW9fvj8IJvpfzcs6/4ZGbdh2hPB
i0bZM6hZOAoDKP0I1J6PcUPTzDOXd/jWbg95CvHC3xwoEmM9sYmKWo56ErI8lJ0b8TNRuobghCq5
cV4Afyos3Ze3/MRnAA4nyKHWu+1HP+i8UWFOmCZ8e2odTF+iAeMB0RXeAH9S66dfJ+MEn5crP+fC
hEQVb+gxYwkxRVtgvws/hTqbhWp5cqp26PRCwkznX4fXqzLXTkXzwCyXztRIO9OuSKpO5vTxTeOR
sGfragBXwyz9DnU8mfoky99Pn1EFK6iOXWUAn9XtsF61SibixE7Cm+aNBWiJuzbEt/1FVSuE3E8C
EbwNKQkLD1ZrcCYwuu+TP8Zb1qaA1J8Z0v9uZiyFot2LK2prB3sOP3h/zkBiVKezE+qYAElMGSXn
qBuSHELorCpz0r6rhSadWcAfGQif7dfSmvoWMj9cxFuJSAocR6bAdICYA/wuNXg82anlNl75Gh7y
U90Yc0cktaKHymb/RjgiXH0qVwbhQ9jo9flKC4hqG+BmV1gH9WXF4NjJTfgzAZCgi0R8llEyJiuC
Dt2965jAfsmqBWDb078UPklOWe/ZlgvxeB0T4pcyHM3MRTixbKtjcPcGb8ylVLBczviEfJ1dZ3Yr
HFsiq3+vsRGZlzA0tj9o7zGLsi9Dccyu/URrn0+u/FZY8yaZGAPSFBweB/4wnmMMvrkyhoVbxVSI
XQLhwdBfH+qRaEPh7tMvTFLRpMsIxFAqp19prvIO1LEwpG0h2DvOEXyXnPcDNl2UcbjKc6LxzZBk
KqCSfV9+lq2PyNxJJWD+vnk3B9WQxi7NrtLf/hSQbnUsquN2HKpCZCgNaDlzOb9wADyDoqKikURF
qJE0duUTh5glJ5ub6Ea9ZP6wp8/1gftDrt/PFIcRl7YSg+TxsbJyaxeLFxf6IGPoSs9/cku6lkyz
92QD4mM7H1YJ+Mc8+zmZ4NDjzu/mKVsuPa8Cy2di+yDMIkZ3o19LFb4hxXdYvw0W/9+uEAOqeGOg
WhKQnW2fuwuNCwRDFbcv4JDi3KDaTYvfH6nZKSdbZwAkHU8iugpLMsdmQQPWXmCgcuHsxLZmhLUm
zdmDwrebtFMKGHZhTJqNFNXW3bJ9IGTc5bWfUMe0u3Nof8zPG+1TGMMWCVaQ0JZhGjPJ6B6Wa1GB
7MIv1Zy1KmG2Q/nbjtJtv2jX4x/eLATaQUVREgkbrDL+QlBulA8ZbfeE80tZZp6mUTRdEuW3ehBg
qNfnH2+nW2IsXdUyuS46uHDtFcgfiJY2p7pZjSm+pMR5oAsrjd9dbhPtk0gTH9Tw5ZrRVPQwe+gz
PmwYicKl4vcXbJX4SmtPU/60OSmzqAUh+1WEUDCEmT1hMI6al8Ma6uVIhb2Rl0ty1VOFKqirV4nn
vVTHkSqV/Blh84Zf+NA6wsVI8ttZpb9WoTvUsFzyWL9+05+W1XdNZLYKqx0UHhL+ZQn4046cvrRU
Z9aQ3NdA+bTP41r15DxIycsJwvkGUWRURGfwB393XM75fu5Wlm+dRXtRrIitMcokrqvo+N64/zPR
W0v8+i/QpylXtVDVon6KvFTKUE2YtgQSF8rLC0asCju0lIftScSLqiFEw+mxOqBPBrWJaYlUOI8p
h9FJS/Mr51uc91ObhyTMQhdGQHqX9/E+VSntNdgORpj6cAsqKZ/l9BDbrpmphe+cD7d9HoPN5N8b
qelk8pQz/uxWT+T0snoIgVgfFGcnd5falOFSXqbf1hBKThuW8q8LXFlen+QICow8BYFW1vIL3Vhq
I1A/ayOWc9ffT6U1rZ15vPURo1/6Qw5JY4L+p6Sj1jBNV/xLJ9DFmfSCXofr8i+uzEu7uWgwqlQ7
9YEpXTukvXEw4Nut5RL3Ip7Qvnx0fHY1sQTfNna840dWIUFA6KV4xVlG3PtmTDS5aQk22v6iBsAE
2uZoKS1GINFuA6QdcENYIqE4Wqb3xmRyYZEez2RSJRnVV7HEvakUY8Rk7fcpkKLugjSIuPIq8BWO
Ul0YPrAXdxjR0gKDkVmNeUnQ1ClgHlS1muFm9NR/xE9KhRmpa6XKhVg75YPDzTKt3HN+otaqx1uX
jPjspOHEXgULwbgcQGhj91mHu+1nxaS5yzgv7bOqFLZCKmTl5PmN3qceqSg+zm1Byzpoct8hjw9+
yujkqTEite2lbc6yLudtObL+5NsWZDKQkIyhbnI6msJULMOoBH9helK/V2zJ/iBk48IirGh7paMX
T+a/rjsJvLVjAXVycgTIAdYZz/VwwCPA+uae5KY6Ue+tg1NwMXKlOF+S69d+4sR52++UTuKobrGL
+xqEzu5vTO7vNgviek92kYo/om9zA7O0d43Ine8+gNoiOMndj7iTU7C2SzqXA7ASg/dQz23mvLRN
vSMd7TwsVGrZiw/77Y3juAKfw0fQTJT1d3XJDZGiurNwLPlWZSz+3vLqSWbgnW/1zgbn2S6+gdgi
tm9GX0+D/WHFJNlJB4SpibuVjokFqldnOQIb3J+Ftl3rI8ZT+uj/3R845EbgyPuix686FIVriwX3
DYDhj12wIiIvlcsbE5BKR/hR4htgnZ9wDF1UdDOWx+HwM8I9QlSHqSRa1ftCxOH0opzjFpHVxbnP
uS2OJIsINFSvY2xRts5VqmJhy9jrBJnkaFdOXYFaSQcWj23qIiUehfWnzJJfFltyXZ00YIR6xqBL
b99jG9J5Wdy0ca6f+DuvALXotwDHyhemLvR0MR08liXrmWQc7LV4KwmuhuVgs0Fej/DSM9QqmiYc
C6blQF9daqj14nwWbYZm80doY3inLsIR2oHwb2uJp8OFUFew4Y/WgOMO9N1CGnRCQby65/T31M2p
WEBPM6R08C6gdv/Pb3Cmbqfs7vKwPMP3N9VCsWVjn1e/xZ4uS1WKLK8eMQvduOKRaIOShbrTaklv
989p+wxVjDqFYaaD1l87+aG8mZWEOSdoqi0wM9rgPjdSveCF+1Duzx3AaZ9/pVOJ/Anz2tD8h1bM
CCFvC5OgOxGiJXBaWYPLv9mY/B8yCQc5G7OHvb2dolNnvk/EMRIN4VJtUfKT3v5uckD659yRTeuo
LY8M73a4Z1ByO2dseeFlGdGrse3BPtf0KUUVH+HSRp0kBM7zxSzQrON6Xkf7vC/5dyrUrOLAQYaz
04xD5FaRasO7ca32yDodJ7atnGTK/QfRsrWfV/9LrJDx7IAVl3xcT+56Gnip+Y6hyeUf6EkZT+ab
6iRwmvjai+SnF7K+G1KdL5uwkSGu4VZnsygyYGrv6EbHmXLRPeht3IlTI8bNSarBFMw+8pfh6xFP
n82lv+nTfUNTnwgpc4fIZNHW5jNLrULn1p5pj4l7xIvsk6hmW77+uejKfNAWRhdhwuCqA//wkv5e
ewbDY3hZtF/3V0pUZtVhvmJVmLM6KiOsocZt1Gd72xBxBuiSvHU48FLn1o7iSVX800UVo4k4vKcu
blOvwxtme0XjyPjh4Fy+FboIBvj2UJ50wDGCXbk+0O1Oqdh6dsS2uIiy7KSiD2+Li0PFLBc+Mhnl
KGxW6h1Az8TqNIdPriGUK9zQTdPUGSLpDAOIY5VkFSpgIogYT58fnMJ5RmZH4e8IP97mHlU/0/3G
KCqkpPapdPA/N3gsMoYXN1TcTZKbQuLNVUvVZhXTndHL2/gm8vmeig6wR+NGdbO5GV/tXkyNwIPP
eRdEhcigZbVs2tRGBjMCF7vS6Q1kRacnXP8eLpFCJA4QXxYv9d7uDZNwEKqqcwR2RnNwetr81EJl
RT31zU6Av42DTIWNB1rAvPD5WEG6imG1H2vOjNeJYYOZdwOeKbwXGFHAYBDbZ1uA2LBQ3XFmgS2H
mqtS5lZwcCi6PuXai/7U+3KF8Aqxpmi2INp3Jh10MeIQgEK/rDoGkAEC6mMSpaFZcfLN45SGm0Xp
Vyu1tRbAkX3lyKlDc5EBjT742Z8SvdxxeKJ0p2C9cciSYaRcyj69seCzIG8cFxYetCctToXZqOq+
9Ynnh/eZGCHM7LTJ3JvX3wjT4LXxMJKM64hNU3c70daElcUbmnRLGIQS9ufWb8V/gx75yW1pi6/O
7cpw6WWnBgBRp6KzBIrodYJx4Sjj7rjznhcLnioi9vH7cw7SUmOboefXMGttSZult7dfN+S22zS1
tPwteQgaJg1c/MCJUlUbWM2g0WEGHcwDTxt6QEQC9Xaaw+yon5XuuAr6Ld5oeNlLHZ9LiyT4zfDI
bNhJHvFahOHWRvmoAXoYErfi1R0qZ8WMxmg/ZVYlXHFlupMXznKPb6GT83e76nH/TTKSWE83P4dV
Sc9RyfGkkfu2W4Escyk99Y81Vqp6xBmwfWD73cBG9goyLLgsxescAsXjCP8OaFsmnr6zlJdE4y72
F0EtsehsJv35PxBA3i1WsXcRpi0y2SVZfQWvmc9UDmin65lVbhuCqzV7e0no6vTw8CS3pMtM+EV0
up5otQDuIBNw1wMV8b64RIXgHo7b3sWamCyXsFw5pTu8j6v1xauEIwpaCVli3p65aex9BueRLYzC
XD5YlNox0gV745yAQa62VmQukG5B4jCDvexJmK7bNt6TS6naKv4VO50hzLD4jAV1LODSvDdOY6Mz
gWju0VcXEKyAE444XRAA6jLoBSpGTGYpJTAwVvN7J+2az7VY2nsAc+o+HvWBke5sbm+qmeAkx7Fg
+YZlWmT3VXnB9RmcanaaWzx8dBmno+pqvZe2Witu+cIkxSDcUL7/K/stzJ/+cDNyQuhl2BdFOJg9
Ipi8PkPvXg0UTRqzGQ2oMWy/MYLZq+YdDaDht7eN9eFo3y9s3T15wrq4iMw170kKu5SHlmPnWJhV
M6W2P71PGF2ZzIjix385fGAOCQaXBmmJU0lhAR9jEzJDzprOmORvHryGP+ewbeM23gQHsoEAgsZJ
KUHpqWtHvC11dmXt6423G26nOjfH6xmWTKvVxQ0Uhcxe6lcqqX0jJW29h9wqTqwknu8vxK3pegXu
PnTbMjGxCCXbi922Gl1TFuEtcUqjv5dhxNSAspIdTHtaaTJcxZHMdgt9ZXbcJDrqRogT1cKYajqA
4ckt0KYEGkW0ps7Na0tA9vmxS5XDt+7QKWTCeqPXrDEHoCMCdgeB0ZuwoOdNVJiIR546uusFIiqc
r/YgIeO7bigPHaXaEUcnNQwZ+mB2kJiKjR686YPQxJ5dCVDSBUdBL4NcAgyjAyWo/bsumvW0cX33
IwItDaQfbn9J++EFfg0oBmaDtXcEsqhCbEZekQglRG9aZpU5ZeT/YGTC3m/8+3sOguczXXvK7E0q
U4OuXA6BMLMGJYh/yLtSEqYzJRIXarvZgkmtJTaQ+BgxYdz/+mc41xbLOhyfZp3IOwOpQirqStxV
ihwp8a5J1QF4xAfFU4gqyBRRwaIc8slZVjAa1DVZiWq/0MnBynXM8L24NAbRklU+2gcrv8adTqFg
plMmrUIhARjv0YP+DaNQrJbnJj8R1cFy2DiBIWqMO/iOlvlc8QHqCyjKaWVoxbLEHvnGaMJGOIXX
V0bbwwEX6caLnfRsNe8KmmcMsNpisVfkVlyGH3IZvkHFCkiJC1kUtG1yk2iC1A4Yn/xLpSwf7wo1
R7/J1ZtZquVncWu+ZMuxye3xj6SJWQ3CPvSqLaxHumJzJXJBfRn5i0+1CksA281HRRg6350H0wqX
MP+h7H6Nu0MJUe+jYhDUX91cgMYiJgqhTvE6dnAZx0JqXHf9Atvx2cC6KJKuaF4z9YnxfF6RLZM4
7XAMyDnkJHnPzq1cmftnvAhugoRb1PmLjlhPt+Uyn2r8RxPnsTRrZ5YdDgB/ibiGfXzbYnQQStXi
TTT9iCjSYojOq+ElBp6ccxIkszQuaGLLJ+B2WsOBVkF2iTZ6DcCXM1FxcIQ0SxdaU7kCBPGz+hW2
l56+krWt2kMuavcqQwPCA6XN7tQXzeRS2sbR1Zde+htY8TLADytHEp0lNLJtafTKPkUvrHwpmenu
gBoVPYYwy0x3P+lWzKuXOdww0TbcWaeDS8RBomS3ADVexkvlobTLe/WuIyM+bssscsgxc5dZpFsf
YjOlVoyjPJt/VHKfMQcT4To7Khr10rNDb4CoaYuGBzirK9GVUCBn8U3nNPHVnLbbv0qtjG9L13G5
SccYD/k4kTNApr3f3AZg6kPUEfWWth8LWGskRuajjdo2+f2V1mc3gbPRv1iC885zy512RWBvNdC6
BpojVyCLtvBcnNX4S26zY8/rtM0LOLKpWuSFg7YTLL1jtkUxSE8uxOiULsKCZQmAHivDlF1R5ZI4
z18IKPr41NvK74wgsC2Kw1VT38RcBC4YxwG7c3vmw6usUcIT6Y3cS5cMd6gxA56lc4ZtQ4bauObg
A9L4ooytSG5hxcHxBU7+ytIPGxsnqcDlsGwWJp/C6KSj3WL9pM+ljmmjC6hKCs0c2nx1DdAPU8ho
fQXVdci+U3qMjgpPUQWZ0lGwLu/GFA2XcO9TLWf9dOeCVlfJnMrsvmiHsaC6tD6kZbY7QQTqOomH
k5Hk9+BEeOXzopXLOxYBsuDii9aZyLjoAn7z1OD52scM8ERbgI6RBX+l6SYpNwkXwx2XFFJBzM6o
yMP/Z0H27QuXDGes4EFbhjuztMrtZbfFK3dToqAS2blEQIfN/B/YX7NdRjkwjN+jF8Po+rcGuKCO
lq9xw09U8ijy80JPeiosd7L4/GPx5qwujQ7waVQEfcaaOYkUCRYHVXLnK+KhPAWBlcCBTSX2eAdG
PjhBBoWwzak3cWxMCAEO9kBeRKzlzOQ9Hjfbi+NU3YW+xajj5gr0KCUI8/FuIoDzmf8jdMHn0Zzy
eBM2tZ5UqSGjAaz/GI9LCg0ND2Soa2lAi0iFGhXERXsX4ksTcowqD5Tr18+HcMkNLih3pHESf0kY
iMeREK+SH6E9F6qFLfxROdHQGvmBD2EUlqGchUbiN4heVna/Beya2qN/2w+NW+xZ+jd/dUTRVWIf
YICfxtbBwIeecRhnUhOzaJH5safeJ+l+0tlBbYDzXeKo/3zESztbCuO0WyLxq8UmtWF2xCMkCKLx
rclG2Qwo3x/puHjq7imAVXfpEuvjtf5SCmaW4BWr6wKxv4Gkf8jG8sm0yXcVnXZkNdSw4lZDXF3L
TzUZVyE8OvDR1OgLdbadCtLVX+l1qytz7cMc2DGJhJeDhAkmm5PvvO+5eCIHudXpZmf+6XPo9wGL
RuykmI+O/FJpHrhcof3141R9KfYpUlgp1WUxWdYltKKtlgklkPZUWk2ZNdkc+a8LdJn0782od8l+
4mqpklKD9G4wIEKk+FHuRawENvixXS47QNp1tbLfGvKi05JUU9CcSrh/dznpPMDda46LTk3tVcge
CauiuLv1CJW/0M84z8U53ECUMYnyy+dmy70bko1Jv05VrbTF/wFpu5vj2Tkv1xmjLrjKuDV5XLDg
B3AODIUgaPEv1cEO4404TjRLcDSjXD0BVI0tgt2WZgLZhZ4seMvG/+E8HFzk5H7NqeIyPrFG+s6I
/yvEV2i5aWkOxj0eq1UIoHbbT9ZhWqpjnPaD/RGfT7wg4UsYkONqP7qvu3Nhyb55ijSz8IKifxbG
YTGjYS/cPIsaR6V2bwATHFW47MrvdSqafcNuidkmRw5jSiiXuYUeDKnG3CJDTVsZqT5Sn72VT68o
Tm2SJT734OUDkCesY0iGyqV67igA8wbVljdrHOnhvgS9HxUlvNXTCxeOV92u/PRAiPDDjVEQH1wX
c7rZrNmlQccelATX+y74A99pBoYY2bcOmpXofabGsy29Ai8cugFKGhfWX9geXD9UEzrYkCoDrCRF
XqF/s7cGXnof6gjSwP/boEdgdxqzSKfiP8FG6Iw/aFpkyV0MMH1DzSXfp6c+jwxdu+KwReVdw+2n
4ozWVGUMIMT7s34pZiSdQ8LvY0QVGnhtwbOLOXcViBKCbW5IOJ6i5X7UVyaZeGN45sXD7euv4x/j
di3wGlglN/4vNXqdWBPQu7vuOC8AT3zosahBYQwtVquQeutif5lUPzOLNF312SMuDaESX4WJWqKZ
Oy12heb3Te/pXbBQrG2RJTGrVzLLEFAt5bJHJ4VVyYj/cs+c7y4VECkshfjlybpip4lG6c7i5kY8
nhDGsRFdd2yjgfdH0iKQbXPAnSw0DqV+z1rJN7aU29IWZOKacwKo29Oc4G4eqruSunaUch0E1SY2
lrZsze+siQ3b1/XumniBbyMqVOoKdyB+SqUhYfdtyLjGOIi9iudO108oOx7CI2r664Zz8zAklRXF
RPndQtSTU0rrdNeBmZUE3CEDQ6W30mDpyBBExrnn037UE7w3DEXRhbIFOnGkQCJoufFVsEGlNoQx
v46hosh8RzW741x2W6Mk35KDzeuOODTBujDGYtnx3uITPrNHWeb+LKvhhy+PBPqYRu5ZKNWAzeJh
JP4rBKc1gth+jkh+LvzDXfzzpVYiZABJ2bXyskESWdTwHrreaW3I2kcg9EWsbYOe7QRyi1Ao6Z70
hpL61RNfwBtcH7hcBYWONaTISfaC0skigQfHDnGaoOLLoUQUfmWStoT4BFXRI2JfJv3GfW34GFKG
XUcMY4/EvNG+tS1IaapsISfwWV6ACDBXsuv5k21BsPnlma3HHOcruBXRNOfZgRTVaE7JL4bnnQPg
W1QidYa+yRkQqCRg/WPMwd8qxmwMs34ZjM75ob+rLKAs1GXtHAduaQG3aIu3x4pnL2tA8R474M5V
lDBoz6wieD/EJkRjROfj2VK3kTnwCxaH+fANJ9t4kRBWrR14qfIqyxBUvH9GEwUAKo1jkxzhJ+LX
DsUdZh7KzJj+6VWBZmnv8X7GHER0zzkoe4afOTHiGzJ+tl6RuiIeV7TvtjPMG+vEY5m8ev/Xoo2u
mhSrY4Dmsn4uDh6FomD3R2+2RaAhkFuFHwizVXNNYuuKDgITHURkhyljQmP68JnKUy8jj5pCl3P3
lAkMkn3ZyuZ3GjDs7xz5sIDGzHFL8zw1dP/oaUNQHdKY7sgh39560dov12eAV7IonO73EuFzsBCE
WjoZhRnLZiLWdTTxepBznLy7IptgOLBlaxSzHTmP5np1CJu8hZa9t5eieiTKdFcL54zqfYu6R2jV
kIGrG/rOASHeedKfhfvoffznlc/w0Jxso8ezYDsGZ4figqgSSv7iEfxAvRouKfbVig3aRoqX5PoW
ij+OYhHgZpjEFuYu5uDF68lndqK8xB9a9/ll0/sKwIw0jj2ZS9xw9rmg9zEq2Io0lBkVWJft5SJM
kYs4keD8AgaI0ZFwB/cN++Q8I9UsA4L8wODgXUOBBXEdwRxvhG706V1aV92HdCN2dwRk5UCb8obH
1vWiFPgEkmM+AzXqoS1DVEnDsvFWWHdEI+2MkBGRRoPzGQasNq04O6xVvuw2hgbNZ0Wnp4wjpyTH
oWmPlc6xryjFr4aTHxKqJKD97ww2/OVNpA5k83ik6oNhdKY+YAAriLH/hwR/C/NhX10WipJcI8pz
iVoaQoJBkeu76/umrZi2LwbAxrgkrV/Mfl5n68Mugzj4qXKVx73svWXnxBYngrTAUZBzr5YeGfza
cCYkJ86ucG195lT4UTIiYwhNcI455LfWKqN9JA3+13RlvbNwYslpitSADkgB+ILXk5LIBavK9cPH
bwaK/S9MuyMykLd00rRbAmImhAg3LhcnzhL/HcG4/Y/Q6I8dZCElh0HSdX2xSagqvO5pbp7kQ/0J
Ttz2MjQ40nqI9kk+rzDM8hxbAauRWGyG5c/Yxc6SzuyMCM2Gnq7ww531vWGspqfHSV4p85g2kuYF
UUwkgpij0jA4+Yc2Pph6/XFj3fMOOeqvreBdWvPCJUS07FLfdnVSXxlCst87gn9p8oOit7lQWWl8
XKyA7wcMR0wvp/5VVPv8+L5kieoHXYC8oOP/6yNWB0sbx5OONez2/oHe2i3gBR9simqJH7t3rqjr
5MosQz3zXj8xwH553fKZzmZNOdq65iqAJQkyupO2ZoJycDqY5HQeMQ7qVkGmzJ14S+5rQlnaGVlj
85uefYxe7eChHK2lyTCyBhza1KuZ+vyMCCJGlCbTxI48T2oVxlJXeLbyfD0JaaTlR/Z5IYiAoe7S
3nXOpryngLt4ihkVn5JHO10D1Yg5t2R4x9OWLFU6Z5k3f92F2AbnPJ7pIO9boeRclo0jdPl4x8OP
AjmKij77cBRv6ZyaOHXR9233z66DvnYtF11V6hg97k+mj5A1nUtonAdGWZsmOefJlGiOC85hJ5wJ
KtuZsRexdC5fjP++8Q1WadeHkQKIoP4rEtdJd5r/XUxMbhn3Pu+riwchI+hzgk6H9pvw9sG5Ngnf
CQRNRa/RCHzLf76LEp006Gm9SpXQxxnYohfGr4HMmTJMyYgLHryiCCsMNUY9Ogl0z0jTFVRumggV
lQXPpiyOldugQkZwzTcLJ+fpBND8IFKwkyXC10bj+x7PYpPYEetQU/MVVwbaLlESFmXEahrROra/
WtUCpUT2iSD9dd8yLXDSlWvtxl4ySsdL4J7jlleKEAgPCyfD/bhM2K7au+deEXARfMxKNs7upmm/
/CNViskBjZbtRk3JZLsqwQwROdQjJxWQWyG7glr7+Pc9yDNr7+TzodzjMT+mD2SztM89aelYxvQU
2LTPmIPV2Ccn4FvI53jnSz0p/W6XCeQiHOI/vJkFFsgx2ABkK6WsDwWXhTzaA5onqL2LqDGXCZOC
RZufu5KMDYEe+FT6VbEz305kIfNT0ip/m1gJ5VMo4CMZOLlVPuQ+61X5UeMTcQ89XC1EFkFAQNgH
hNI8Fe+/BZV2PQ6cvYdolr+gCRXsZ9PkhIF6MnmZJs0htLC/Wyn2enfV0oogU4v5IXISKJCb5sO3
4Pii+wupnn4HRYFpw9owZ2leRe3ASDaRYYu1oVPihjQKlUsKqS8uJ2FLVaUvZK4sAf4PLGrAmCga
94rEy6PeBSL6fKajLJQO8UEO2ctKMNU+Gvcro6JkHVz7T+SZ57Knpt/pvoGCx6/EAw1rSm4akdo2
Yw0XJJ6btU8Mi1ol9pD5athavyxYz5xXBagNCgllmWbN9v5ZMpPxBWO2I+5yJDZxf7O1/8KGECIi
AEpgu4wqgQ8mtb2GQDE7MHGpSHyxQ+Uv6j4Rr9xoxWEkr5AawNf69rl7BWFs1Il7yaacPTz6BNVg
58QwlKD0ZpRMDmUQpuelDGUmw4dkm2oTHla3RuRZMNBCZfMycE/sewmTmh7jbdf7JJRKWYEaMeX1
D0zJthkv5+zIT/R5EhsHNcmmeWEimrld9Gf9xrmRQCzw/9MAzTgmPZCD9IBRH4Y6isD6vvZTOz2P
/QJJ1ZpgUwIfVRiu/w0AOBG9Eda7IJKs31VF+1GtaBBlblrasPfUKETqnREjXi9Ypg+x+y6aeFa/
RPnrmnn/EMWv4ssPDfZ5R6nLBFnN8lkFPoQVXoFQp8gBY+Zvh8q9lah40NQ0x+pckkgMd773Enbh
Nwu1z5vC5plM6SdhGvEjoRKl8i79oM6kXUfjkSAlYXiYyF5f5iJwaKtzxkbfebRuuDuWr/ZXgmxH
B1s3dcO7Oydk54IKdYXuLw0eoVvaCRTwxYxHZCNqGlJp5R8mblcbJXpW7PR090gg27fEz1XTm8QF
yrPK74Onxwy4vi02VH2HT4g2MJnhzx8KwUjgeJI5A6u7B08IT4F99Byq92j8li35V5yGZMZGYdMy
XxpXwz/qkbolcdjrYYZte+gpMCzUB+B0uM0fDmprMWXVSpWhdGpxFvaEz8pdEINemMoLk6VKqhU9
poC4q0XgU+Bml7u6Oax13fnjVu0Ja7RRnAyb75kA8esLQbLEalM3C0aopThaJYi2ZEUT7nNsheJ3
DoDczML6dlcEMcePX35ZWRJknwp2ZTZzCkWQpVSEKGnrAuRZzWBZfB0iPdzpIGR6z9XQtkHTryD9
c9LBPsLKcYjK5VGJfOUFN9XPvME2a7jK6dKo4hTRjtceknPwlT9WJ6rNFEz0VZu44Ui9ETPybSOU
efjSaWjJJIBSLBjG22vlTY9NUizFdWy4R5t+KWFjhWVlBDNNomfKGkX9clN4rwULCbCQqmG5pvKg
S4jdXpj5e1IYTWlRPC/ddrEqOMDYNBmO21Etvdn5ANosOrRfCTpmdJQySV1Ho0KWSxREAiWvuEUr
lP74hPQGvYqmjS3JaT37TjIOmfF+rBOQPaWDKVALAfHU+ldu4QPf6iiBtIhPG4VFsRR/V7+JPItP
+m9xjQ8ZzVg7E/BCT7Qs3CUI9Fj4W9W/QBGwZ5tHqpV7MGajJ3RvNk4PiUW7ATr4l2u/7ZtyxNOA
lUBZV9BMPn5Wz5sA4sl2nueBBSpIfoXA0F0OSTJ/YYjr4B9bv49tMjq43xsuDGJF6HXTM6pA8oWL
k2dgfZKnYAMDhwddU3NJyJeH8InLL8xSPzj6ro/oUtg2a+v7hlAlMOFlrvF4UjARg9EEbb9z75sB
gWMC7zTTRm8aTDEZlLLuyzd+lSOt0rRrL7XxgHA1QwzLNgIc27TS5fY1XaybP91Kvl42CDbzqRbj
faSakg635h6eEaU7uhBd/ENXeKFJVVG5uO0VnXuOTt6TBreXbUavkWQGBUQvCk7PWxcdtYG4zCUv
UKB6/BkUhba7dQF4h3fKjfm+1vf4IlCtmCla1mBjmp3vnPD2Qm4HKodZXxu3lhTTyt0YQWpvYD1j
tQFlNsRj+MyxzOW/FffZJBqpL7qzEwWTPqWTvFdjO85mXd9ZoorcPtHG96qUIYKXkPMZImD5vqzX
NSwLil5/qftoJUWRNsBsxmXTWLUXa4XQZl9U0GneXZ/w+H6nSPlumeblHIEg2tjD346Vyq7zJ03L
iDRAVq1cn5zW63QRHC0oVAmb6Sy3lmVibZjhpoSaQwEC7EMJbnCDEV7iPdxL1NIuZxK/oaEaCJjy
ssnA6K/TQlmd9hdgKt9EyOGbSB7VUsDDNX2szXd5vB3SvfP875T2mg0FbGkV1gJU7HdSEz1CviXJ
z15avcie7UI9BxvDvMmu0u1doUTrFjUo4R4mZSROqGDqFHYywkwzDWCASMdx0K9WlNbF+PPg60bf
kPRZKWNi9GD/J7cCG+rfRhPHVd4/q0gUdm7qQv6nYY/n90WSIEulcRSBt5hu6CCiobqvR/LxiceS
ddNOh+PScoYTfcEM8XHG2dY2EPwi/c+ZU0ctZds40V3PnfGaY8ijCWwmIcF9i8uzhW6/6//TUCyN
G6Q+t6WtiiK/BmZjC1emo6MAC2Etd1OuvCawuluIswHL8v4eHgIHLJRlXUTVPh72mZh95KJmW+3k
8N+0aUYRkIOmYytyPqXSZInY/sB9QIk5vX/dRjmWBldgdlE4narCxh9HFL6Da8nalt5rasTYBw6q
TB7Wqq8pFD57EFBLmgu4YcFfuqyIZKVzegKJ2N8qyNGEQx38aF4Uw3IFvuPU3I6ghI4Kn+feJAvR
KijcveuQcxzTmmWJUMdpLOyJSNGnwH1zkk6ic4oi8qADR9GT2WFHp6e8w4kNXQdmk7DOyFUuS9Xi
B96YWogK6N7B47nNAXdhuFDI0Gpuq92ArR37qaHyhXJY01N432i0gfXrMGWw8tGx6GnjD5gkJTl0
KA+iR2dkgeZw7rpaYAgAnXiHwcyj312k2FInnnK51H3LAIzHyTKDHkIn4g0OeVgPdCDno60SO380
ZGmHVaU5adt3LgbMA7NQ8AYabgQC2fzyAI6BIlJiLmg2muObxB9s4CgHz9IpQ1Jm5neKf/2IUDMn
2lW5NJ+Kz2yzfwxUS0QjpCWi8MKgYKZkDsOqGlRF7WOG3eewse3vIB+bYtcwnLrNQGNLt0EmSyDA
zgBI0lb0UGpSktPSnx50BhcR4kIjPgYtUeuySj3JvweCvIGSHZb0oR8yJx1jqGSskeH0Z+NX9hhk
HDRP4a3mfkjWtSkf26X7LmDJ63ZTc2eE8i5CaArPjM6Z1lzL6ZsD6hHfKiTa8bkq5BWi/07VX8nj
h5YPLLyqf2kUS5aPeOZ6LJCgG7OmrU4Uk7WNXU8NIf55WSxIlXyBQ0kQXfLShyMOom8TUT7JYKvS
DkeConVN83K2PsdDqvQd54axIQRRMgZ5CZgT26w06MMqnUelMt5+QeZ/VNV0/DN2EBF9+plQYJN8
wy6bRRkPcqErHAojOEy9k44i3y/MSNEKIio3xR7pqWRHwU3VtQVMVMQvlpB0IluK3nU9VbFwTgPd
afw+z+sKzhNH9K53O3n9hxheOTFKDvLZ2nZRVN/oN8SazvGVC9/eyFEHLBhH8h0qR5GuBljiqdUg
Jw4CvxpHnSHxNUSdYY/DxkUNHsA497Z6VJJ/sAtBilk1gLuJtOlOx8HOuvUoerPj1y4v8gfD0LDd
sTNOVJOmwGvC0PFwR39d0jMyoIaESUfeQCke9KAd1nu9kJZE9ZmzIrXnKS3/ftlC+8C76d6nAtIx
ivv2GNZJbh1cbJ/kOkZHL4q6U4DLFbOepAgEoUS+DLDZqTbl/vlnbCZhFfNcY0btIBcxtewtbZpi
WjAyC+cp7o26MvvXMlCLxXBTBUyFQg/Zx4ByWhG299Ri/XgzYp7t9XBeXV9vG5sLgRG8LGC9cLrY
BFSLVLM2E9dd5hWypY+ni0sqRGSscu4C5am1HHeKiopcryUVVMcc/PwmmZDrY6HWyqzx/qE7o2Gv
i5/IO1LLjuiLlOTPa9zDZyjS1+NjDKeNIkIh15aJ3ieT6ryd1fdQeqZMlcFXuCo0CttpFjnw1qdB
UYqytX4kvEcMVYTk7irIyUEkSTAFnsEJAhU8+NKQu7v3RbYzK61+J/1jQMOwlCr627YDgttGUt91
HFgVjF7swG5LeGXUqlm/Rb7CNFhG74PyL8rvMZtbyAp27Eerq4AhYa9HwpGSsnPKe7q3JARvDFac
6PVIeB25tMcr+EuI2WgsEnoQsMwzcKHxbAe9jmnRbMXs0OJYcKtPK5VPO7KR2E6bndZG+SIc9Shz
hpzCYqHWU4+GHfeyAwg00Z4Wx9pnWwxjrp8oKUJeBywc07ipKuDz6iMTQA7r+DAQ+Qo+2bqrCG0g
JRhD/grt21GheFXyrN6wK3rVvrhxnEKaG3I2h/txxnuD11bg5DEbGXlr7nCi3axAJjZ2IHFjRaF8
SotL+xQTsdnwS8+lJRyhH6KwCV/MekUcnecEzV28N+0fzAxolxJFZXi3BcP0wp1A2tmf5Sq389M8
Om7cbfuvc0e5szJJMnwyD+r1xD6ZT9hRYU55ttxp1dgNiR5UEqRIR0bHztAvEzCkWuReXQ6mn8k3
EerMUtsuvra34lSTZVvQy1unxFN89/yJQtM/9wuFCnNPwgli+qlcpTPPrnhOsdLYUpj1yw4bpmhh
2T8bqvt432swWPOZXA06vG0hgGDMz7u/cHWEocZsU0ppbI+qAFEgnOalzwcGIKZrIdXGzAjyxk7E
Fx9du70rR/fBuIHi2AQFSE28YmCJzy7DIFH+X7fX3kiSwKlGrPC4ud27MArbtyO/cZ1yWtLwPkth
Rs64QRRknKnxMUtRZbRH0LEpVEJXvhXfT9S9mqKsCl8mfLoXPHk6acUtjneWT4ch+sZaOp+w5zp/
/3OaUG/DsIIS3vSz+jaL0bKMvcw62w6UUnoIcHK5BZTo/bwFIFwUe89aGUlZuiinE6CvXJV3ct3h
WDOtpMDhDRtToP+sONol2QV1hthUVM6dGQJBNOWQmhvh/lPJC5D16kD/PhZov+K+7m1LXvR1xGqK
Fbe8S7iaMj046gxZ+v2Lf7P29/wljZlh+m6HppmZPqvrJKzNYj7Rcq0nzMh27yFLaGveR3tCuyen
1ufl/zfTnmFIVNej97vdeEJawDsyy9/PJpoRVv2ZdZCCkkEojJmT6y3qJoRMWPEQ+raKkYuAKDRa
6fxUjteO5upY/s9ZeGSm2kjm87BeOPibtyQHfvQ/7JRtlgmP2r0MdxmO2VQhGuW3vYicldYlTzfh
uheZm84qhm9JOqOkMZW5BQeDYHxueg7/oPn8cNRHf2jnQSv0QqL117FlhHE8kbQtqMcIJH88sCZt
49gIm2+6iVI95UHa7uYTCIL9tokdYFcun2jfvLN83XJcp1BSvIAIA1HPLRlG1ieRCa+kIz/ZD4vB
Ff8DuYwOnvsXdiCyqjTErV9VOTxWEM3oRSX5e1f7A52C42jh5L/QhT1aFi/jBQGiSE6tLO9Sp9Jk
ZFGyZoEKb1ljyTCVoAi4uRzt5Z6iGP+PN03R5aQLCj7wapK4qPNbexE3hojH9NHlUYTqXO/GMEZq
DvwXTzYopAiILxnZpghdpy4NC7c0VpZSQRM5JQ18Tw0q3qb8fnBQ1NIfp25PkBTY0zsjNcL3Ls5p
v0Sygx2CLjCXEHxQXQDB1ZPBSS8v/YBaZj1gvJrSKhW9XbQG067sus13ZoR65SlKzrs+PCwOE6kZ
wnpVF6lweCZKGwgMnAslaPiUfHOr/pL56I+0GYTrcLK3QoK8Jg4ja7XSHqxeXvsQaduWfzvsAsqN
AOuRY1tarp/5Y/MTXKSK9ek/+Fwky7JAdGVgzIIuD66Nd0d5013EgAN5KevfYT2Zh1VaqIu6SGgb
I6O4ewcv3QN247TbJRAdgwvBRSQiCRR+MtwWf/vpFAuOfJh6tZ+rpDiRHxjcUqzhQNV/U5f0FuUa
XxtM+vPZl8h9WMEjZWdTGXFBX8v0F+zvgvwZiI/A8bDuz4/wkGOeqd6rFuXqypHPIbiOpNHS/n8J
PLE1tkHm4708MFYNaV6wTIub0X8ChgJvQ+1wNsZoXSaKQ3YMj8qLygnYxktet6ueXWlexD4I7OfR
VPRX0w5UYfKH+PzwRRBe2C24p/bO+5y7RwwhSpfS1D+CiawUBcWVI0VPQqEmT4ORfOEKufJhQWMY
om7Gskel3/g6DwqccsSB72DB69T5uvQ7L3D4tgtywXinCNMzB9+txi6VIWLrDj+kOAz5si7zEdzA
zxZxWpCjN8f1pdVXiwv+bYk7jdaErgpVbSdOu5RfgPTIJPZ8aohkXUxK0t5Hsk72RFQAnYyfAEoa
/cLM1kO/2p1SXEGAD7lRElPMgdmhvdn1GfrVTVTx0/BGMrHXO1sqTPY1b6NeqhVzKTnXTRW/KPas
nvDt6x1nHdpGxF8EF93pnqQ2OT8If+Qz2TkMceW5251KcLqZmO5uq+arMVroMqXMcTujvNRB36gN
ILEPWgv7e4kN80TVA2LwE0R9Ce6vniVw6og4IWlGN1oumFXtv+JAIQYm+1xoEOI+Ghkbc7/QmG7C
FgkBwcM71w8JsbTFtB3yxA/e0bIdb2Jhu3DEt/MxScyUSEVWVH9Lf3FJkwlI/cgRTtOLdSLr856U
BQQfzula0kNvb8IDTGvbmzM7IRezxUNGMf41PKKJmIwxZ2X5kg8ngNv3Tcu2nSdTnjF2idCiEc74
vt/XUmavNubjsCYat6+yJ+s44nLtwyOK6nq6eKIFp+XjAg99ThkYWknyc2NTtg+7YNy6mLP5YuDM
gfbGwl4y5BwcAiryukwPZIjq6d9OLRQIlvv4Irg8vJKAvuMoArdzF3wFvKtJ3nayBrYg1PVIb/1t
1FwiqrrL8L+xC+4bK5YGqwdM3MbT39uzS3HT82wdsB+SgJX7z+gzTRb99MFCnVBEIitAFlMI7z1J
NBKoOR9Eiy6hrisgCCQimBsH+A54qTGJ22gHtyQycSRb4fGgaw6QdNtwYKVY5u5AZ4irBcVM0Typ
WZGBGvT812OFcZpaKy0aIdSSAhZUt4Bv3YGI4EaMvEPa/li9KbNBu0X+9BLCMU6x8f+1FcHd1TBK
8UpH8VBWHXj/Iqu5FcQq0h641THRZk69LsEQiy4wQrCW4jS1RYPRoA01YJRqNGd/UTD3XV/oioFZ
TeAHD2fHZ3yaCJ4dWXv4y2+yq/J4be8Q4uEYIOek0Ddm8nIUKMyHEsEE2nSWfdn6GC5KXEK/nLO0
yldJ41yXyG3QaZ5RlDzukYb0dwpafBfadWZqgktOtIwnbip5ufZh8SDk7PR++/DzlnPpJQPhz4Tg
JcEpPz9kcCEQbL3wnNhLn93X5NFA4sJWshGP90qihZVlYJilnnU8Hr3D9ApjtKdV0Vxm+sfmKiyi
TzOdxiLdDEe0WEAAH9gH4zD5jUCToRqSqDQY7xwY4/8i6VNScUb60GaWxoafdKXBLM9vQIjv/uio
VQTzFcBWlsvii9gYIyKDzlodN76O0kGbGPKt34UNw5N3k1EXYllGhFSjhLK+/1/rn5SFXKZ1vQu7
MkmRmf0Cb3YPua0uGBP8FWhwMVMKylmAsg7YxkqZXePbcoUlY00OWXE8lN4+ZcY16Yz3ncCsw5RQ
GdzVcKmH7ISWq/MJQF8gZY6/2ZaMB7VSrlMuoy7LugxxtchamNYIoWawBnbUFBt4g3d8u3hknANy
+ayjqgXtKMIviP+6yDGdVP042phnVloRneyvFp4snkhzuxTCA7mCPklEWNNF03sXVY6eDQyQ1Wzq
JxaioM0PI1jeXT3b8h9635KQKXdVNkvfahBvEgDasiYOq6IT43UFf165iG/DBFQ5hLkMxB1EqMzs
nB2X7HFAOe5EW8CImw+T++Y2a1R6oX3x4Sz5SC/Nnq39xmJGxxm1AsFnqRpfD8ByJ8issvXI+zTd
HsMOtAthgwvDtQG4vCYZCcSDOUIifaixs+qk7IuVJkNol4Q+Pvi8OE7PDjvN5DwRZhCb/Hr0XVX+
5RJCTAULb+mVZWwzE+1WHcbqy7qbCBirhPJ1+3whymzlzbFWvrKIJV7HAeop7JDtZvEn7N9/piQE
uCfn34IAhszU8r7qVI30W8eO/WUprlHkDtcuYrUgHva/NZ29G4DOYIn07/P1O3V/Qma/VdP/rLsF
FdOimvZLEXXuBebJZhiPP2kyZP40s7xQeHQyI2eSSfSe86vMP7VXkgAm8gooEBPAZHcJC6bmtW+6
BmrX8BF2+vhC6R+jLNe0Krz5q+Ys7OefqL+ASLfXjG9k5TU0IAELcj7869FVzghOLK31VH7Jvlpa
xXjrI/vJVHC1aVF7aE8fzFyrKhKXXRcaR4XUmvt0RK8R+Ml54V4q93GorM+IBSJsJSRjCwqDpRFR
BYdDLvPhYYCCuMdkOACegFQ5efJXdyL7ZqdH1uL49LLZlKufyzmEXGwSH1PrEOELAiBOrmdXJEz/
jpeEDr13lg7zZDzzjkhbKXLxeYZXkXIZOBs4wFEtHnTFBYKEwENT2FW1wByVEH8zGT+c9N0BU1lj
XXz8mZfaZ9eJz1Bzu5f9ANj/KOzyi8DF0e5d5j+zgR4NmZTd4tT1OVkL2uI/Mn/sula/NpirtDhp
ju2QNMAwW7tgGKjddxKFHhQyz8uOvHh/8EjOjSXy29tXrhC4Y5uSU2SRw1ARreHlshn5myRMu4gi
lt1YhSfiILCpaXk0L9RMZtUAJwblPYLsrFmYefMZ9E1A44Nj9W5rmH2CIGHWg9kOhHB/mOQEGiEp
qyYIcuo+xrdbUaN0CsUaQBFSTyIQ8VSAGNblQcADv6LYd1fu2RHuiPV/zG/enqIyU3O2BdVp+cOT
ZuoIUiJ5d26+mk+7O++4yB5qQxeq0sNpFPzE5FK/NJQ9y8IDtAayC3peQ0O9fBpWWPNNflKLJm4I
LBSGNNPfgYD0y7OI07uqHcbJR2akKI8gqrNxC+It9TkgusYxng9ZT9p6mq74/0/f/ZT8L3gGbiaQ
qdx16A4taoda6XqnnvAmBQd76KJCKZYokLcniTjNMnBmzQNnG/93PLeU8tNAq058kCOQ2G6YtVRw
dNjqqp6CvdSSJc4VjIvcUlMRj8WoXD4mTorJahgfSGEEwE83jW4/7ksWIpv5tBOsXprt8VLjXSux
0NprpPwf/sgigK8Hzz/0y23WqiK1YfWTj4hO3eYrCtHiG5dbEk/ejayQm6jHFU4e3QDnoJ6xZYrG
v8geRjyFOzVsqpwvEiCWoTgjsjLvNDyjNRBXT173WuB8RGHn81CvO9l64h/tPTB8d7/lsZ70yk8e
r8Mwpq7qNX3Wd63PW8V4orwGuKV5bvXA13v6apKXNtD2yRlRKi6a7z0+nzTyU53tozx37g4JvmFh
I5KfwqI9ckGX9gbOx97KOG0v/fq95c3mcCmRR5cM/uTNUsvyTnoGOH3mYQB6gUpvga6QJ/+f0zp8
MPI3tXwHUpL1BuXoFjERiIcaURm+iXZpRnnQ/O8+dj4bSpJrDzlf5nNKmICb8Va1CtCwizZHByB2
h1fiIV93ng/TQGtLYDWgtxkaNj+H36fy+xJxqFTWy6hkPquY6ok7mgHrGf9cjvJ9vlmx63hM49lP
EZCOf9a/brnVDDWtcPnM/+Uc2M+DMQuEdat5ulxKDrRZd6zIxzkJeL+5T4nWMMMDS7DnaM7yBEvX
c93nuP+VMwFOZgJixQciCiWOP4BpjVXZprK9dd4p1MN64MN/ZyzMqm3ZX8kNdul83IKnHfxN/IZl
vknwctQqPPZWTWcvn2kdln4jKJ/x/MikBMFKJ2PMf9CtEP2vd/j4GJ5i3Viy+lRnDSudOJm5yFgv
MhHhHnS3cRrLiLysu4EjSrPNTHQHXt7tjO+nOmwCuEAzqr4rrIM9PrMTs0y7O5hnze5D/0mUfXGp
rAgxbl1UsvI58FTOnhKJuTwRtDb5T8j5cSgZ+iEcIJXLDS+3FJUzDdwx5SjXKmiKD4D/wrQdu3Vs
mCOzMeQJgnyEFJr4e+Q5UpJdKo2GX84BnsHEQsYNJksF+DebHZFBhLV8EpscAbpHgD+TKZtY/VZN
hQxNK1BBtAaQCqA4RLEpOUJ6Qx2lU1WP9MoYLRcNnNtt0xYGLzKltwdsYuZkt1PU/CwV9cLZVPtK
edJsDy8Z98xrZGcfIG6q6RQLHEvBovJdBCM0m1eIf8gGc5ckS8UXNElNaxLLEIyCI5uAbQwUzqB1
OEPoc/+zu9JhXosCbnlawrgcUz/nqstuPZ/YbL77Ry3jXMMkU3cF5saP0jUBqu7aMq1++0DX4cJy
G34QnFC9565/5reF8kBzKM/3Z520RgiggUW2jOVKpGL8aFhSl3S67pudE7nNLVWBkQSJxuTPbB8u
CgWOE8pthe4gvvl5cydx6KF0sWk8w9AxrutQp5Z2dshvWgJSNgk6mQgxSPnBGQaIy5K+zWoDv21Y
fFrnl0FMCA5ouZ0fl8zv9SCK3lIcQSjYavR91a1gxMo8C/cc2NynHKEHgfWbSdAleY5UrFllp2Jm
kbzJdO09ZNU2p/hDXXov11Tzv2soyQ8eyM+g8974XcX2YiSGkKoNAAGRZ1JHEPQ30EiAqvUNKft+
dSB4JTZKdF7lrKP2lG25DoiDnAT+kYjgrgPLfzFL6Oyc8hNIzguTUGQwS+yJ9YIe7Mi1miW7EiIc
S0fue1I6vHObuL4Ryy0/JJqsrvpg6CF+711DSB+wYP9uPD7f74MGbDZsuh1qWpLy0zQ50tXYTsbs
gzGqr4ufkwDqzcaBx4zfE7GYZBdY6zGvEOBNLF/cKZATzYaQ5LuuotVQpy3rWYs5QFL7TkbMzL8h
MD5Tk76ZxOu1gWqL2zgLtGIdnPRaUa0eko15spnC0ynskKxCOKRBos29dvQC15Tra/2Vg6K9xcY8
zxpE/NrVcIk1GdB2cWDnac5zPaiF+uTGSS5vxdag1esHKrXeXRLcsUuTDgi3q8PcDmgyrEVIy5eA
7MCk2lKcJId+G47vgKMZsSIMfUnA+HMYUtp9SUW2gJzcMXxdIvp6Zp2tJ8hvYPjN/fWLxLo4b/GJ
zuiqONjxOByig5ecqFQRMRDI+JGygRnTXBl9EA1y2c5Hh2bX+eR2feEocOyD9fIFfrLiTdC/QjY3
7MvVY/FoT5+JFo0+nvKmWbFnnKKW5jBpshpDF66NNrfUJjm65YwHxqpGWo2uJ1ftAJL2Wj3RSvOZ
a2usZ9F4QxrV3ms2VLxoVvx7y1Vr/mrFm4K9XJ9UJhm5RGDCCplyABhtla1xY+8dFW3P6q42nmuu
urCQSJMmz/JfqAHUBoeYEvCLItygfg8O0Y8GlFWcHC6SKWukliv2ig2RkwA+NEeKBNg8hXtB+S6i
qXqcLhiVhiLA7GcvcSKOsjiUe8BTbX04CtEUKBQqQFIJx+xoK3Q2XdyxkQblfdvjrxW6r27KneOI
cbrvRxle35sabNec0kjIoatVNu6DPbBNfdIUUdNMFVQrhgIM6Eewb1XmESMfz89o/cb24Eisvo1k
6WndHVYnzY0Nw05fSCFIK5tKpCFq+pNvGuv+QBTSLrPyLgJcu9V22e2OgJ9cRVqarHPFEoOpRXf3
75g+xlGTufWJ0dNf3gzItzs/WSyWGY9tkjYcK1yzUoH2yuJnPyYPhS0eFBXUzKESIm2WtFI0kEP5
cSA6X+a3IHTIvQqNkiTC0KnTsIMaeM8XWFvonePFCBWLhox0wOWBlZPwsc4cihzVqjg0jzGyPA3k
WkkW15cM5uxF6okOGUTzK6es4H/DdvDIhqAXMjhtelL3mZPkDM3vBoAs/zWWSxv7c5+9gzE6xTnL
+E7vihRDO6pYzd2mSL83RTbpOMQzWw3tqs/TLq+HPqnc536It+q4gNF7U7vZzfOXOTM2UOyySeE3
dH2UyVLSHob3FHpBBiNqRfW4Aj5gM2bc94o77BGquYvsm9MFOkoeecuIWeYd9KKLDnThNbL7RLBY
pRWCTwiloQJ76Hbo95C8ReU26gGDR6bxcpehvOPTCzsyYNAjY0YG3v117PtSefj+5u/ZZfG16e9H
BeAlV0FReBHZGpeY3Le5CD/5FTv4cRCg5JzRmZyC4GDipbjauTe0RiDL++mkvonZr0LUHHWrz/lD
JU/3VLSlnC4hHmDE9xoQuGyTLInj6SPmdxOoWBZuLu5dI0HfUlG22bIAJdgEzDymyHO77dBSPcF/
nq4hZ7MdUqgTTFTOReK/9N6Co32yrPsIxT+vnuB482L+kGczxuBsBwUhXMd1MIW63NuiiBt+Wpar
B+1GEtLFzK8JeNxSY3jod3N07pfFD9SOt5CuO2ksdRk/drUw2JdcybBT/7JS/vVTF69wp94btb9d
KC77gTeVbjEUJ/+mwXKQ9LkTurrmmY8G2pasX6w4nKKy1l+U3mVY4Ybm3tHdM1E9lXrLoStpyaTf
ziuP90cmzeKzOSVvML6j8P6WAHSifFTrBqHWWV93xnDLifiTEvPxNeifhGadY/sYEoV3WVvT6Gv8
s6y9es/fEmt21sDrkwC0IWA1IpukWNZsNjp5VWibVQy+hss7P1YfbpmIJBoRHHBWhBsf79TpqsDI
etVTwRSqgGQt/5/GwV60dYYAdOXgfBqqzYWbmB8apzrtEdzlSa5Y1oZf/shxPZrpYBgLAf8NcD8e
Sv6Q3gJ4EBC2dPRWvwtatFVsUAnWMk8yQZAq2b1hF4FgWo73PGDn8PmIZfrz2h1ummXlta9dtH5s
IPJh8DAXWi1sXAXruCsOeP0pt+/7k+dmtsXcF1DiaYdKMzE864ELybIUXiT7l+ykQmFO2UAvHrei
edfwNg2O+meomnlDqnhpZbRc+aliyjWIqFYgxgwgfidSh3YLqhTZXmDbAF2D2uXCskfk8bVLGfPS
J/nLZxrczyDaKLYMY21/SVJ56X2ohfr97Rcm9crZIrm1cmy+97AKnDHW+z490ZmUwX/YaQLKeSBL
0Tq39q44duWCBxXG6Lja/BdfnoXE25q+mLKm/db8Fg/HFDJiTZ+HvrQGzU7EtoOWXlfplDsakVjK
eHE04gwbsAbDEkCsULHFzf3j4fKGMg/dndFhCeXlEhZ9E+ibD4x9V/0Ur0SivHOuykXVZi5dHXqo
KUxp8fC9KxJCeO0ncNQFZel6VgEUU+kCE4USegJeYHjH8hdX4OjRSivAIn0FMDKoC+rekKt8CTM7
sHmB1ZFM8Rx7K3nhBmNDG1smORwJ/+xCum6x2QwE6rPebIR3cqGlCmxW7ApOOWexBLKmjDL0oxBW
V6oMFstAmPyCwKEh6eLqBRMc1hq0rjyvOOPfOolOWr1wK1TLmK3NtyoqiRaOVdHrPkbOBGHesDOu
3lJaNq9ZNfyTYYkduUG7fbSjtYUlt3hEsNtN6UKytl6KSXE4NJOPsfYK+mGZSa/pSiD4woAubZTS
VuEwnAZPQwtO5JgYJEoGDIaB0noEPeHLaVM4rEPFVyJ0uxUBsi+cK/+1BwVAkoNx8xQ6D6h4dbNb
8dV/grDqdJ4/jKWA1VPndMxDJUlZoFyDy5j7i/5tbAylLWCn0aPWjVdUTfGbARM537wb8l4603R7
uPal2ux82z1ciBBbJlTFcdoTHifR2DzFPDl010wcA9Yo4UGFiCyRrCWyYpnHAslYYSfbmsaa0rGK
fs8BeKE9OSfKv6SvS7MeJnLNLcLuYTQ1PdPuwLDrcembLwKXHdocLP/NXpoJ3PBT7bC842TwM6L7
/BSbwcBCPKmcXeQtRqAg4AMCSWdIti6nktAL454AbJY3jYx8Pv9xD9EMzmJXwiOI/HzBxOAxk52E
DoJ8X5Y9h0uqMqMyc0DsRc0So5x+VoUH5WIxHF2WP2lpIKpmAzLSDVSR1hbn+0k0dFKZlLdVnfpn
/duUupZ5kzX006O3BevU1+lDRx6RogcR5UtcxIasg6KC16k+jacL/bj5YJVoVRPIBPWHYIVgZLdd
4tCRn1fiB1+W/tQsaBd5+XuLiF4Mhgg9296OIcHhFi1jq/vv0kHJgEvZqIoeIQ5DuGWN+YNeJ3Gx
i6UgKlwDU6uHWpXikXk0bPwWGf6/Sj8iCZn3demMk60SlTAa3xX5ViHu4cg7c+aphuWM99jkS2gX
2zi+OERQRsqEzIN0qQmUDrMk23OEtSmHSAJ/uaG3C0NyiQpJwDxFht/LUtDv/2shwpkNCgeGhr9u
uKBqu6vsbe/d6m3B55J7kc6ltSa/mxldMMZ2V6CkY2dGw3zyMxSu/Kda6wHqb6RI5gowek+MkQd/
ouoBxJhZZyExNoID0y69G0A/KKT5uSqW90ENPyw/OY9c0iZS1JxUKDW0e7dddo6iR+VzpTF13oQT
UydhTIHvmNf540TmiaU/eN9JJgJVHcLOkj9UNRtyqtyCVCl0kps+lAiFdkRy0i7lZPqec1H21Uuz
3wN6FpN/EqpxWNYgAyJHMvi24ulW6PhTh+SWumNMSTuJf6qdFMGeYsGX5S/3vN4IU03YOL9rVBDq
FOCIGsr4X0DaKhwIh5Uq2UnPDjf3zy7orFTuwOVUVcciyvTfUfx+RhmBlsLyHNWptk1uM8REjk2+
5NmfWhIPXxmxxKXd8zolpifT/7tm0bPABNtGzsRkXsmjfIghOH+7f8ynplPeWoFlGsVQelIf4C+N
stNmbCOuZ+MV9cchV/bP+oXoS4OKnwLsk9L9kTGjV9BREhlLmIsqYcigdYMvffGYPyeDQKZCOZkV
TFuO5cNzVoMvF5oHmulH8bBZCWH5dzyNQ2Sz4DJfSJk2m1uYeFCp2Lsl+Nal7nKIi0tmiRa5HwAE
H1bjN9mZgYlNzssfqtK0JIWvMlaqPIJLjj08jhazDWWIeCWP2XhITcClEgMfp98Ogl3d0qXkrKdJ
bUv1z/TTEI8y++YlLZn2zI5kHlM4xQZ1H0YNHAnwis2BTW2hFcqxeaY9BrCONrO4lS1T75RuTZuW
F71CFThe8dIYOZrIxCIgC/YBKzEousuHLkqEuNL2Dnit/NFkjB2q1jo76l4IAJPkcG/jbwW/w1uj
cGCLibFBkbZjpSEbEoMuiTbHzcRNLc846CZ21EIGaKM+Iuck2wMqXUcCoajdgSctN+zyumIR29OU
9eoZorToLTCga++KNWhtRAiD1oKaud/rwTvwqQNxPZDbuq5SvPECTbdomrI8QbN/VnbCJgxJ5gyN
ByfPEOwXnRAgztmPFKR/Wa2CEdLfqcV/ydq+7XODnXmLW1AnaF78hq0mDP7knfrlmeONBEHz8wwH
7SuxNoVq7o8wyiv1UaYVrIfcjSYWn16U5dBVnQUQbwMhNY69RMmOWu7Uy1GQSN6MgZ2wZzZEkg3g
V3Eft91OzkqxtK/ivOSUFNIgjhCvaCnLIfAp0o6ZvCdRtVGyDPmVL+DBUwB8vLeLUpgV4SUifr5c
7rm03bp/d6lTmanB1X1HymP8RaE34TFN7ogNCtRR0ZMmr0go9cMUu5EAeMV4JK3nC6IknA4LtpzK
dw3DgCLcKvLMHJSqbzdvl3MmOHztuF2ybpnXk1PBh3q8xJ7apV9cc07WmPHV6uewItZsJW0/0zSI
OGte4M9waLTPuCBvXnCHUvgj1VyDf4gR+F+EhczHkAVheYt3Cm85hyw/8d5aP0J5SmoKcp6S8kbk
cvmE4XWL/dhpZS2qEcIkJkcJyRKSsaYUZpKo1Cbs7ZvVDPk9C0GFvUzvgMCh+/cNbqJvhLLoDwIq
kqaK+/YdF8lKrKzyt7bqcHFpBOX2k11BSJZ4igIz7e1yBLP9fMpjwjjGwLcLIOuL1N5/9UZNolEp
QFMQn7XgfATKx6PstxSIfLdcCD7dNT7h0t1jA3UC3UynDu+kYpcLuYZmsvQoRn4CIt7gVl6eyXUE
TMXVEwVShSmf/TIFGOxNC2hbVUt1pidJpXmbwM554LUkqeMFN7g+DsGXsuoGpkAFI2hHJeqfbq7J
/JbNWM7WSup6R+hi+RskWTLU37Q4pop5HMtLj0Kj+1NOaP5Erpnxxg7WyXKK92Ge4Mlmh6OLJq3V
OOw02FLfhu3KtRsdwyzn3NlktCnTqdmTBT0NELtedgUx9WtPf6jrNQdBQ5UdfE/J1KlkYZyLJOlg
ZqnBP/ykP9/tEHDzb5DII13K7rS2dJSigojjjHnuwbO4ZeibiMWYpoQBUW3Ea03RhLGUCxQB3u+N
g24cVL/3VB+mpeU8PUWnt2fDHzfBrg9khtSIw7Vt5LasDEMKNv3DbXrlpmTBQtnopcSZe/wOflBk
ZfdcL/UfRh/cV8OmjXC9bfroxCKbWklrN8EeoV/Elt9HC8EQuhRgp3SQjqbmUx5Pu2o6wEq1Mi+m
AFCQE1ekRC53EcMWSQhcipvGReRHBOouxmrGu1j2kRo7WGitKPMFki+R3cXmBvVHkp/YRJ5Klh3A
w9NRDTptkvYPBnJfYpt7a1ZysYmuP/XusW87hieylg3CIokHgvJZuaLmM1Mjhu7lDmA2Sgh8MuZd
i1QIaaUdXXEk6tlC2guwru5qTRt9Rz89g0qcjekx25xCFZ5Qj45Du2fPCSLnfN/7BdrLuAHQDyem
ovst/A03wLsLNT+MZMbKaDQ0MsTyKcYOPHqyHfVPp/ZwADqHG8BZbUJBZwFK/uEFXOqFII7ugr1y
i7Gv2Zql0EZK8AX0BOTmqQLOXxU1Sd1mrEXExHhtgdGdJPENErfd9vgpbcieX7A1vSvJCtax2sOq
X47lX3QdS03qhH3UnXV1nnqJQwF99PThjMEYGAogEo0gC7TI3H5YRuvUdadUKaDsuGrDEFUHsJVu
zgneyvmNw5XAWOaKmunMcLYeF9lhi7ej377J2DrwLRTUi3hoK8ybkILWO+AmfyQLd1yWWwrDKX50
wzw6RXIdtxlKN42HysZFehU+m41Jq3rp/DYpsHF0LePoYO806V8gpJGtQaD5IqCP/V18IwKNIyEK
qcrLpADylA7CSkBtzwSWxnlDuTUwkcXmVR3/dCHt6eelPIlPmUvGxpDOtCAyfAspy9npbjXv2ZPw
KH3ZW5v0G1Cp8P52u0AygQFxd7JyljFyE9W9fn/e+rWn+dvUo8h/vDcK9BqMQMB9BT7fhV28E4CL
Stx2u+lpLfX61OueDCfownhXRhTsTtgIf7MGIS9VAk+T0yRtg4yEwfbLsVfQkHybE+yEiMt6et2g
3ZnP3Af0tvxAQKscQci61Egz2v+o2gFM6MI3XQ9DnVYwn3dKnXh3FrmK3LPb85alfnoYcZ5qmPC/
6ac7MSJniBhmraKAz0M4JPsJajCsjnuBEe2zp/IR6yrOuCSTuqErK+L0NIlcM5nkospkWPsG04lh
y6d1ZFhC1lHgved4mh7Cx8uAnLcHmMmHXbxQPg6QJmbGOyAl1l4omPkpiBuoK1csx6MCvIGmwWwp
EyGO2mtykVmg2Gba2tRznEktKSapSQ+N7CGM3vOpdscsD3Y6a9wGC00ZlRAKQvj5A2migG5Eero2
vPRnVuMg6KStujMAmuP5PBU/+AZ8/WDTTHCFAJeOI+ZjD35MF7IRehTwu+JTdOMcfYvrR23nImzF
97SkAWlKC21pe7Rr0PKhbPzRYADrrIlQHCg5o1/EkwSxKRNh0EQklquq4xuMMWTik/okepWx4Sp4
LX69EOUeKj9kKEmtygd7chasv5vII8FrlbrTEaHUj2Mime07JugVkNQOcdLB9CqE2kAV3+cT8hI0
/XjEwxRhfYXQEiSyd6buKs5mtR94iHN26j9FfmCTwmRgINyJu3BWTbB5ebJXDzkmaiNju7J1xxqD
vwdh+5Z1+X7uMImR58ALj/nRaBhMJynl6NH1a06RkV5jGwB393rH0Cb2tjBoA8+pZ2zCTJh7mqrV
V8QOxE5FJkcdHzWPX4r20kMz2HGNe2Y3nk+7wSwp1P5p7JrqRadH2p9m2rss3PR/8eMYMQQ72B5D
+YvL0ZDsjGcpahBY3mQKWwkIVLMOEHGvWC0L9+ErIOgMhpOE2kLbJJILArS4211A9wNFa4IQogYo
rXY8O7oMi8NWNiHQMpa2BHC5boGBTnL3a+atASx87JPEA4/zm6sdVLRvp7/M9KOqNM8p2KyMs5gH
zu3JE1zh8IciJ4gNbrJSYq9Xu4Juhpgb0D3E5zceoNcg12E2Jan1uxUqQMZA8ik66tBHkRxkXmPB
bY3gUBmSX+MrNinJJLvj3yM1IDql4UMcF+3JsnGM1AX+SICqrV1Frmp6NcMMpYsOXXJzeGcSsgkC
9Uo49vOnpmXPcr/WCqoSLTJ59QCyiPLBzGBO+J4vF+uLK/qis3fnqRKOTZmDGuMBANSNTOPm5Ci9
Cnopig6FQFGf4zs3oVjlUFVFomHI0rBTQSYx51SLiVCqZdQ1dSldThfsWmz1lhSq7iG9xmoyY4St
4Aat8qhstju21xO9/SdzfqfCBErdSof81Uo2xaiGTN5RYvGTTTBmQj05dmLQLrsDg25PEbwvD7LY
nJSOY8F12abzgxYErc+aqW5lyad607pvZVJ/1uRLRQ8RLtz0czwaRBQqazuFRYdDOReTDumk9H9C
dVBtZVWZnJF+R5WCd9AscAlQn9I0AzfcaTqOlLliNuU1UCD+qADfMBuA/5v1mV669Tx1e2SZWk/r
b1TahQFariE5EuEdKec4wa6XvMHu/aTOwdjDcdEYEMKHYvTyP6dT+nU9dTJ65pgc4/SsTfB0ytf2
c7nsT7KqNKVOQTDP+UiVNF6xR7e1azQTnWYyhq/YcuT2669HZ8+Tx76ikfq48DYmr0m02E+79Kxx
UtlUdODrHg0GpJZgz3q+2KX2oHlb7mNbvTDGiBJCHpa0+sajupAupCejC+f62rKxTnJTz3eqLi+r
fLcHFsjmDcmfF2FgYqdL/iu4YCMslw16smeROIWlwAyOz7Cs4BM3aAu3YHZ2laaX9N4M+8NXXhe1
lutFmHRNoxaFrXL/4BsQHteIpcVwLAGP/02jXOXiQOhN3sLBjHLOoD44BOkB4+C8LvGqmifzBnCP
JQQHX4O6LF8QKn4+X0ftXCXnmQVG1GkrMSzzV/8LCs1fczkPoK4y7YJGEmmmgAdznqVaoWKZMdQQ
unfK4d+KyVFq17G/2yAsisUM/B6f/lf7fHok8yLiE4nEAqvD8EuCVx4muLojPPeToJ9fvAytSMqM
9iGP41s6VojKNU2XMklDRQK5cIQiR8Gd0oRqqVXWorhR9bpwd3fektxyvTekI+3SZ29Pr0OyVNRQ
17hl18sRd53O7u9zYp05hUFA1bDCdvLuEeiLtioYdlYGpgBtkLID53YvVW1JAV6jEozajptIWHHy
JGVca2LOyxJsTRgevQSwtSZcNo2L6jv0cNtRREgoPSDABL2dC8BrQSZzjhgkThW998tQ8EhfKnoi
A4NcD/cdF4c5LVkM6CJ9rBq9DGbjTXaAjEX8BQoZbuFXc4C9tKPSX3BHBHNgBZAoSxShmqcVQlyn
y76IH8tQwWdCPc535NqzrGZn/bNJWoMbnBCtnushq0X03hS5PjfK7FhhkBytkt3MybgLn9LH3ViR
D8iPXOCyOVFRRz0iztGPcJhMdNVEtu0Q1dTtLBr1+rSN1lWfLkjnk3/+xjo+FKg+p1n1ATDDvRNl
vueKn6RBPM/TP+yKOMatJcf4840Wz4iF6J0l+PJUN/SXvBihV7EvgGzEdW/JBcs7I59v/4nFe4Pz
gOvrEyiFS1Lze1bJDbsJsVrsTmwqq87WerPx9uaXI2j6Hb8pODQVrmeVNwAVfxACX4iKmNxRZbz+
fM4MfSvZRbnGk1ePyEpcamG0Je6Lb1TW0tev4gggE3Ga6JpbH720Ni2Kvrn4M5j6uVcKwITINKR0
plNzuJ+prXjXpZ3SEYwQgZJTjEIH7YSsYm0Abtw7+E2//tuuTHBCNciDGb6J6pGD9YmMcJPyZdSz
HuizSew5bHZzsz6IiByAQPY0WoUXa1eb22KSs0bjh2dJtHjc7R0lA4wBQfnx9hRd/GEFvDVwtwSc
7mvNM8UXMrSn/dok+1zxgvxnMvdw19iAmA2k3SYCfpBPCUF6iFgDWGxvwzNyqE6pOvzNLusLNFu9
C5AaxDtMlQCpyi2/lvzvZEhRmXsAcpZbVl0XhV7KXtMxH8L5Z8JnKpcQdnPzIvjfcW0w7mlA2T7b
i+Vi/DZlvIYybk6vPoZQdJ5FnFrunV0mMyIhwDqRiAJo675gAwXEy+rYsVYYJ78VjsgjKPFK6eLh
Va40Bau4n0xILIK3oG42Ctnc8H3WM2MYWgsRhgsurJ+FMZGHBQ/BF9W19kcwne5/qNY6jGJFl2oU
Gbb86KDsYMAZB00GQYk3fQXw83t1AbjUocE5NYtc4nwLcYyQuOKsvk1Bh0l8+cO4ynvbdFe1o/8t
XGTGZHJ/GU7DChFrh6ucia72cYnLnrwTGWksxKLUElv10oYFMktSgMWmTIGclZclJCIfJ/8lT24H
+1wXbWeimNRdDzMdyZqG41365NgMQN/1sxMSaTz00pjnQfv4PVerG7LWwFELeRVe2VcXTYmLe6e+
PVazNqL3+Mie+CPqipfYOd67uOzNCCChAdRo/z7CTPu7XdlpPbzjWK+RZgrAZ4WKGt23m9T89Xl2
velCDr5kj3RvnzGeMcXjw4wm5EfkMpYb3MH2v/VoV1lNPRmBcsFZQtLrW7aasc4WbeZYXMv9pWqp
ogEJAyznuHmPtawDqnkLPzU4PS1/72NxNuIgvs8Z/YAZgUPN2MJoYn/F3PdtEjh0imYBgUtiXMCg
f4UxDcipyx+DnAqkX/k6XfMDKXPs7PXDHeY4R08Ku4ZtMGPBPdtvB7UG60XtRZmG0t5fwebkpS0Z
2JuRDmLTQBxnyJbWb4V/gkdVy04mnLdfw/iU53hmod1+VMa4ps+ynW7OfOvbQnGcGCjNgk7N1Q8C
HUw35hV4FQ9Ki6Ps3dec5q1+fgf9NAO/vREvmxxQ2TQZAvfVD5yeChnRCWuvPnAisZvRHojoxZ+U
1ArZTTUWY5Z4I8lh1ZIA8Kq+mRo49xn96htzZKDeu5YsRvPVcqfT8mmS8jdw9nC3ZGA23AghAu/L
AuBwiStJnHURvSoKTG735DbEqgWaO1hgHGdW7Ph5kHfsUFFoQ6YPRnAHgpbWhJBbVPgAR8EFkDLV
LroNtEtfOSb6pPrcc+bZOetlEOt3bwG+cHlwJA2ulUiBHJyYdyUJDL7IKJIJQPcbKdT9MF3gwnxN
zrF5XBQ/jkOvWm9ttSLOllZ5aDgL4EVPsjucWNUAD674/xjhnICr4GhP9jug9MpoKUGiy2gWZNGV
xHs8ueLfNYPaLndVSiKAZPcN15zXSb+g1eR5rvgXGVbaO5Gsv33kEdjBFRKmkuXWHAzNp9BREC4+
SUGOp7J46je6NhsasqPdJRlu9XcWnIHJlLwavwXUDQh4hcFAwTOEmLy3xU3mzrcvehGOKdF1I+H6
bhitktIoFFfK9LE/VzH6IdlrPx8unDe/txiWsjG9qD1iuhHsk5hVcanATJApFdDfhux1TJFjuDM8
t4/z7UYzuwNwqwC/xQPJJn6O6XCvyF7FielQB05LCkvMVD81OXRXQt2kXIbMyCHoR1pfuKIDVDDb
/Sp1hKS8EU8dDk3ahlD8VqRAkvZ9LvicXtDdhs83J57MYvD7smGj4rywOGwkKEzrfmNAWdFWDk0P
SIWR6MScdQAyItdugsJCdpnPme/gbPBwup5rdTa301+jDGOMaXiGA6uqQQZjfUfoA8reD6jXSPH1
qmG2rQJrbiAQM7VGTWDWgMV3WCpWuc2zbstqBoDzeSxA6SIBCJdDj5BzrYrvS/AxUQsIo6NSV1vq
t6lOP8XPlPjLgEsVTd5mzh+qCCvpbJ2jH8d8O0+WKnsv+RMTTf3ZjY6uSe09BSJY8Ag7DnWCR+D1
MSOvqnIYMrL4Q9tvjfWMTcFZNHwwjB/PvdTivko5zYPowv0bUXfSs1kYXpjwIymf5AKckWUEIGLk
pqhoyjN2svSTYeNqUFRNtylCz2cpLfNQkBS/4Hafk2fQpbeySxn+D7WB5Hf8vjTEv0R9pTRESwRx
l6ppAhyw4xIFLyI8H23fAXmo456uJ499NC6Q8f4yeceGZxV7sUZoFDBY0u/FnfcVCqrloSrBEUN5
awqbZIi1vcBCYh7ZiyTmMC7f7CJkfpNG+lWWNo0m53UQSgV/0xV+ZicFZP1udYAmlEfZd+OiQ0fo
eY46ZtDmVXEtsG2ewhOMGkPrqYoMsgi154TDsKaQDp5GS722Jw0waXeM94liwyVDPvCIO2/MxTiz
85wJBflWRbXQRuPN+klT77c8PUO5onGs8OJ0U3D55E3O6lbwqWxSVuIfA4J5j8IX74WptGsCLQRT
wcSLrKD3GwW4RR3lglsTPEcLOIdW7NGeU/J1mCxpFfB/FY2Ye1SKW0MwVzFhACm1Ds4/jWe2MWUH
1Pr+GTgxHbz8+pQ/CtjdxZqJiFNwxxsVbfdEKmQpDPxf0+gcsyiaNLY6bG2Jt19As9JBdUYRxtwS
phtMwwNMV8hiFudtlzOCfS3EeCf+nTQ+ZXHkHuT8uAJVJiiYepZLWxlyqyffOHvRRcVUx1n2WAR4
hTaMbiRib7E5mRqSgoJ94EF3G4Hj3otjogYEcDWIaW5yW+bGWnTBhRnrQpd1wnEFlVpkYf+qkZLU
FBT6RixQ7mjb0e2vZFCwk4FMJcNHXnVdVQ0ycR0tlaaisZ8/xCdiMnAfpv0fBIJvlUKtYYkE0rPV
gO3yfCG1BlkpcOSU+sKQKw3P8L/RIqDaqEXIqIdtXS3puqJ6PiOOC1LLexlbgSzKQBZXOhfio9V9
f0jKkmYRn8FnC5jyJoppFokFbW4P3egQrA1ZALIiyvUq+6aNEbbalOb2oqsOoowJFIj0NrXKJDgR
97zgDL3VCddTLSI5pygPDZz7Qu5kAOp1MFk4IrIWl/6Vvx4d2aVydqa8xKNReuaNVPK+7TuFR359
O78kOjpsmlj8BmdBjP+LXuPbyjec268MO3QDJnEnYwtRiieENtQBwvJnYOPFN2Kt8ZgVd3RdJYvq
L0M0Mgh6Xrx+nK4GlT9+QmFtwLUopb5BspWYMjIFyGY/hzblQMNTyVBsTZ/qpV95oj6gZhYI4XPD
/N7Mf79IIjWNU5yIj4iXeyU8vrmX8Rh4MW0O5T3UyB7s3jtSnW3PWjdjfvSmV3GnuXTeYMxcoKvC
n2U9Tc9v2uuHDTENucHydnVbrIot5lQw7vCJBzELNIscdD0WyN+SWqPfJhVZmwG1esfqeLqwIsZ2
NmpCPh10AGNwDxEqzS7zl/xP3NWIBqTnSQst0MS+4I1jn72ztzFQhj24u/tPGDCkzmAsdbgVeoct
xHdrQB5LLNk3U+QHs9ROjie7pts7wl/DijguAsEvSNxQrrcFugaIHkOqrYo+cE5q7VTJhMG2BEL3
yB6IWWFIoiumA2oTeHxjDznYZezDirTx3d6CsWFQ+UNUZG0dhuunP54a3XCHDR99WSV2YgujGVPr
vujZYV6s2lTAuNm/wFepVTyHpWsVotSP6AOA0zWUSHgFKetK6frzBOlllLozRNbJQ7onO8J7Y6r6
eSUQyYCPiYW3mc9K/PLJdPjaXGiRCAPZQWCIo6zWZ2/yK1pCuRrtm4ioMm7Hb6S2Kg5IcIXLzAKI
pLiTLwMqNEMQgUS6n0lO6h5+Vk8I6niMG5jCbs+tyapn+3LHrA0Deetz6zLSRCDGJ8AP3F0CbgEF
/qjYMOVHmf/0vs5TS6w3xH+odN/G8gO5pOl+d93jkifugL0BP/8W4gleB+DV6G7euyaTBTE/dSZS
dbwAzdVvejdzbze+say+E0vuy7nptCLbeQ6V2OlNEdu5VLJuXmowEFd2WMFvvmvXznyp9g+Fs+v1
4cLfQkKrLP/46Xiv8qrkaGE2UT1UL8U8dUXKvLAz1j1IpZ5Wik4pOvrhgIFrUY4wAOgAQCufNmoU
RJwNcUlfLn66AloaLh8n5qh8VaVLrW4jIH9XV9eZ5ususzzLQG2RBVxdjqR+UhSMjEYt7AZswGjZ
I8OReLGXOxrY7Ukolleo1nFkPEQde08UNhoSjeRhyImirwsBH+KxAOs1l06C4waYtHTBHgrRsWB7
zl3iHP+c8xT66qW7uCdFaOfT5Uj1UuRP+dSDqy3TLfjPdb4LH29N5C0vQuFdOmbvDCU2lNBqDU7M
lYnaZZzYPRgqXHYziQwPf3vYAZNHGFX2Q4dX0bOlNNhfH1MprlRRv26N4mO6Bxd1O+NzrnaIog2m
VoxhjUKFn9LzX7TR6nMno3y9wmk9sOM6g5Atw6zHzf+2zbFnWrlovCiSNFiCm0h65WhDeW+ItLnn
jWLH2FCyDVo0E7im24/mBdiux8MYYShEG9LRN82dY4CwDegAI0CCXlnuJS2v5VnzJX43JBHD5ASl
1JTnJR2er3dYJzziTSYkT4bKEMSkPE4LeA2U7zbGf8w49ew4NZusGv+Mmqdj0AAxAEUXxAlMwi1A
F5dAD6fqcB4yHjlGnljMwQ0eU7FOsdyGvVQF40WsKWY4L4lAG3Xqp6u1L0gVNxclsR8wJUEw5g68
ls5TBjgwiY6yJK2xqwQ8UXX0RkyNQ2o1KQwgHpqPurXOSZfYeA2SewNN3O4mabz8opqC64N4sgG+
0mIltCLnDvepVF4Bi6XZCoCGCSnVn2VH9dLHP77PVoR+MaYc/kmr6jdqNiTSGzig+ViY9OQ+QgT6
CIFCfSrocEecfUePoiEve2O08kzr3a+5m1JN3RJCrXuRovSRqWWweg2p1SZvdO0kROGO/EX+QL4s
0aKwLyn0GY9ZflIxJTDsYFPC6zMWYzN5O4LQlIYo0Al/BhoEAKIvR6rJM+vBa/4Hvo7b4Mu7oa5a
Pdz4/hSRXqoYmOm1Za7uIkIF1S0gTMwLOzxeYFdUsRaW+f7wYd0wISmZTZaZgI3zFXCHR/XuDLpG
JZ/WtikMBN0swmVFgy2I3A7iEcmMuPtN4Hnjzi7Cz8F9ldE459GydwZ1KVNLxkJO9D/A39fJX6Nm
vZ7lw78No4nCuFMjL3xYVfqyBR8vn4TewxXrqu/96x+GZgeCMiIVhBTVibFzDhIfo3yH99jldSOj
SPQXi/ytgUqSLAAsjWZGPSThfVbJFut2U8vd5armmroqIU7jjg28V4IVFeDn8wLLpR0sCv1rgtjL
M/sMJoopkYPIjckN+3o8Gv97m4nmdID9Eo6Ah/9WoHTZZE8+Gj4E5u7XSjUMNR7MRE9D8iCA3acJ
Prg+6F1du5FzazVeJjpCnxFtcbhUyJaLgqJmSkIaRHY+1ZF2WsVKmLfzf6wqQQVJXVfcJBYjBGTs
Uu2r1eTDlr+TUjupKGGqpnhwtj0bd4Rt1nEyMc98GnpAsSYNhcmzqmFafywiXHl19i75D9fGndEN
0FsTHbLZhHRQ9bh2Bdi3MYPX/7frR5SeTWUC/FYb+JMe8afxfI5GgKtmGj8uk5UI9JFFtP4nq6lb
3fkVspDCc3frHwWWoIiJoJ7U1BMC4KBXgqTNyv7OyD2+DprMEd1uPESgs7Mt0+XFjwxvX7W5L3VC
Pj/JGGJizX+fYxv3QAv9s9gZLsj1kSj5FWA8rAVaQIRZWtbc45tdGr72+dI+w37I93tRqK1/hot1
1SB2aSYDtxtC1PeMvL253zYUCAMm0qTKGYfeXg5aJZBTbDrf5DU1x7Y+kPVl+uZnS5txcZvYma4L
DPd/nF6KQfYwQB0XBvVNnWlo/H9unOYiz6do/UEKtrY/e2dHfY/nr5ytv/1yMomNUJ8HbADA7hma
5ZprZEQ0DFVto4A8wqC4Q1Tz1Iz65Gl24nNzJ46ONZEGSMbnmSJhnNwjRTy9pEoTsGIn8WjWDFOd
AczmD+YbelXioELj3wEaNaVm910Li7GvUxRbuyYeGXZqGiEUtIRG9nvp51WiUpR1Ptfx7H7Nh+ee
jO5jY+5G3Mry7CZ0ZLZiTKxlIu939pRBaofuIDS/79Z30VGaxtqou6zhYHmTWEaw45G9JcXTQtdm
kdWXSNQ/TUmncMIm/bVHVr+pb6QqPEFUm69GMYprH++aKt/ysFdKVGKwhK10sP94G/ZcnM+U6MOo
A+xZgMVNnzR/L/PrGFOi1TgF5s8ms1lV9Ze/kNvZ4Bm197W8/N7+0fyFLIulMEpobr21pjprnTXW
U1tEONOKB04cho2mjF7z/cNbAdMk21q1FNK/1XF88Q4zkE7/DS5/f2nf9M3Qi2lowykZE3XXI0u8
JvwjU5BKcCJ6AAfsewsS8wy7zkyj8OUjgN8TQiaKA2wHjVmPvLyGR3D3oDXEcjCjqmcUdEVYCbKz
HkpwzuCKUpHcs8m7oB8WX34V6dgTCETbY3Tct26F8EpP5lSNg7SBnI1U+tsBGWM+jKQsOZQKcSF+
Dhq4KG5J9Xx+9BB0uE/dvqQmGT9qgZk5lb++a7/ZCtN5w4KPdF7P39UsWeSw1mwMDIeO3VCHRxl4
8L4MNW3FFX6Ru3VYhkBUhnYTeiPZvW/yhM0Ku4MvOnTOf8KjpD4b5LMvvBoHi6lwbdX157jIJRll
gVRIRGx6jtw7/eYV695ml5XsWRpOdgf0gfhvZCUWhjX/J0yVHJLPpLF1FZHs26gszpITuHAWD1KT
Z9yus5sz3k+AU4FJdcNQOfy81qmnJ3K4y8c7gOlvYHMYbwNE9yni97tCTVre17XKvtXhULaEbGno
4nYoaihi+yzYKnszNXjZ0/WdCSOnYB5DRALpb8dJx0WRlWIOXPdAeqlGFz9Ng78aZsws4djJ0vja
+LUwemm9xX7WahTKiEUe+HWP2ILcta8JBGVntNy2H0w5AliGE7kEHM6PBuqgaYDFepGqt1WfmDlf
++krzN7L3KBal9Uf0yIHm92qFdcNNmx0Gp2y91rjz+wcNSuY/gpB90jqhFHf7tzG/AZHxyHHOd+I
GrTRyDgMw/e/SOTp0oVkYaOZ+CB7PWXSp74ku/bkASW2IuK8nCnJmqhHFj6TVCuIJ3E2lyD51bDi
sGJ1cOd0fAicW2Py3bP6n4e8xnD4tyrCMqQL6FK37IISdzlgiBIwMGiKskplFkj4z6GegHJ59UjD
NAHfNxH4MX4UOVCj/ys5+pxJmUG+cVLaCGBhjEwtThx5rDURBXvSW72N16LzX7aWY4/w05IYgwyW
KMusAfjCB2dDcx8roOF7YobvbLLxr8f0aB5pkQ/5scuLTi7821ynesDSuBYCspmWoW4ejfLyt93I
3EFCP66u3psrORTjjXaES+KaYdShcEzxlTJkDQ66I4j9SqGfv4YwDs9FUm9WsB6cr4japsijBBFZ
sdv2TFMy8jKutKm75GodJ9PkcUFutbzbydroES3n0h5TIjs/Q83WTXTchHVhdn0WrNE+wwovoMNY
K9MTgx2upjAOS102mC++13bxv4YteSC8Fr1PSEqXGyQUbqmvatMnEEcXMn00B/xgWc3+EDqz2hF4
pR7JctC0V1X17Zn70GuDMjA0xDgTrMIuWiqlpu1zrj3uqz8cJssCgCBnep39dvjUsdaAzrAJ9Lrq
2Fq+fCQh+txuxO4PaHNDGb0VGskO1vmKSiUrES+gLcr4TD1BsXhBi4UzVx6eimaSA9mTU8ia6/B/
6Uob8gSVfu90lbWQUC8EjDhIuHWsoExrmeiZb/LrHaRkb3jYHdjYzvWGNbP8/m4t4Y8gdLSxLpe7
irRDu0Txv/RLplCyPwi8ai4aWjBhhCwha0f1XAwh3NsTltB3eCwyv2F5O8CQDi7s/gCMaNWclqHo
QrQY9fCOzrfdGTiRj0qnouZAEmZOc8uITy3x9QO2kyA5Aw3diQqfhXfw4BAXnaMCluMum3z4YhHR
/06dZ9cwJ8Di3odIQmGCw+RCgvVLqowJIvmIrjcCVH3tzvi4jaT0OfYikdeehtjQ6tKOJJC/xc8j
9o/zrw3cF2ul1nGujfwQSkqLsCj0fkZVeZEOFfK2s/f0RhBhltJonUjBVflEbfjJJyrVFCw733JX
MoUJNkx8l+RpAwJRqZNj8/qOhHYpYGYIQKkkUszHMAV/uAS28kb2tiKvREpxlQOuuAkVrX4FE2Lq
18Hm/v+QRQLGjblT45Z7MR09K+XvkFYg+AIU0mJFxliHEoAF4kOtqCPSugUrW50FJ58RcdQ8SBLo
eCI32csd+T9d4Cnnbn5lNUXJaCZ3lp2pkuv7CdiYbPeleh9jgJ66B3Wbt+DpMrxv4br3Cs1gk893
vxZKxmdZLHHbWnuciWnsbqG+JxMjQoPjAO56LeRKBVGC6DHP3IECTbVOi3F/O8NUlz+4ddWbZpnx
GaFE/29CMdOOKJyiR4CehdAxNIrllhwD0WzycnJYhBJ68y88khOSn6/hyEZzDYCuJi5xqMrbZra6
DEQTFjoAzLhfRx/30qQUL7AFo6N4LGeAATKfr+3svUFImwnQ6iXYB572TFQi9CK+aBrS/ddEIcXv
2Vu7glk188sAO2CSBKGKi/l2l8LW3OCaVKxIY5JEQRVkcUAASF8BTal4RsWIE83pVdEbi/D+yDcl
vyVxslYJXvqaFaMjPM82IhwBwhbI2mMaUE+qDLrhfthzoYmKzsEuxfXJQ8OOkbR3ilRv6pTfJGMR
o2OVPeS6G9sSMum0Bl4+YL4vwABztNbAkDOYWVht4BNXEG7eiT9LRBhAz8K2A9KRRM4/6b//THJg
iDRAb79hG5vizJF8CpBKVjQGPzo88fF3C2Y/k/xSwnJT1oHW87pQmzaRyOtSfuq1lWIfZOpWgOdI
XqsF8c7PnHn2gOJEStGxih+zQ0TfRVJvWQSAp3f4MH3LtNul6Hu9vERV3tEChjzD8rNeBAE/2M+8
uA51MbOt7M8tMSYvjwY05CvKcw8eLIW9OF1Jaaj519qftpZg6QHQNWKhr3ngBPrMbeOePmASpJrs
P6NgZ7NiTmKVNqXfn94BHbQwgCeGWe+kJu/W1iwhmoU0/kEUd3KKCRJpRkbKBK/QMZf+lngFvHpd
k1TqmDfLrEg0zMr7dDvbcH2zTwfsdOuZxq10G2KksUOeflihK2CYI21iCc+sG/y3zOQVgw0mHalX
nrWn95UrE/oiywsDgn4fLTeSRn5/d1uZfXVgztQnFxJiDtZ9QVzHv76j+hovb7in+rcRpJfpev2g
Airi3uh8A6MZCHPot6NRAs5gPQAHIBGy9CIWnn14MctDT3C8THkMASMubXtPGkUHvw9mE/yjF5dq
2eDWsVInEzWi8iiNMPe7rj9Tv866gNuiBshveCpS3wGoWb7OtJIL0BPDV12TPpANDvJA3kD8cZe6
AFJx94GPnvdi7AYfwkY0YMKYx+OEyAqv2P0ILQ74s6zq8yTmPLUY4+YpAK1UWKFcgUowf8top0jO
517WE9eCDU1o0WP5ZuQhCn+FxHG2EF/F4u8wqOuOE3O51fEc8PTGQnwB9CCOTJFMDk3VtvBJEq63
rPA1i9DgB/WO8m6sSZiIOEEuzy3O3szqe48HHdvbvg1L+5q55P2sEzrDbCiRAHpCyOdQQM9XisZd
uebwNSI5mD+utI32YMHdUan+aa4GstaIqRWPyexyKMyQVN3g7IswvHDLAVpfk6cQzT2Kb4ecK8JN
3WbRUkNmcXd7Bx+8eL4MjM44YJ/zMBCqKOfPRpFC709umL0K8sYMoeSCg7D21Dlwg3McnoP40xr5
zbvuX5Pgb8drbw7yo3atLOUp0KYcjBhFi/Mtc8pVjy7+Uj53I+PTjYDhnJxz7KcLQW/FBdfjUXNS
B3grm2Zzy2DJqVz3VP3LcG6KJdeH3Ajt96PwTSdGunvLPLkiU6AIuhzVVB9BmLnGW03ERWS6/LZ5
xK0lf3mUs3VKux/WDOEt4Hx0NWsto6ItsTAOeSD88W5835O71SHOelagwq8/SJP7lNCqt6zoMkz9
X6u74+WDODjI84e8rXvilOR3SOROJb48363/c1xjbvE26cGg3wQEhsUPFJxg2C8/zf/NS3SDQFMN
Z/bombbGzv6p8nyCsho/rvKIFI7tVdfFvuBVMWRN5zppv7ltt7lp8HIY2/reS2MCoxwq3Ii/mSxo
o3i1wj0RHjeAz/3BThrX8vONR/VNlIqhtyjgqk9nxh1QcHIHRwM1szgIbNepGfHk7N4UfE7HE2qQ
yuZ4KL0C3hnLztUCO0nn+qGWwoL8eUl3D6o8s0iOJqEtIuiefQ7V/q5yO4ColjBYpEGmiN9NVEKm
6E+pkH8DUCGzIABNFwr3KBvZJmoGQ3qaK9E6Rx7q2HjjLKR73LO2d/kJlXC3IZmqwlJvKSJ/Lhql
r4Lk+DvDWkApH4FIqNCqJFCZEaJZse1boG2p8+7v466s1WZGv6mTzFsTy1wPmIobr8iO0LgL5DET
Ks6bNGfP505oHaBc5HcKdMCQ6nResW4sJmVAHHJsQJKpaJOHBYp1FOwTUwjFOqPI9dKjko33JT9s
LTginG5wUztbE9bfyWtqyc8gpcT67fSFhula51NLYgt0n9zAsXMfISmBbeInaPA0O0S4XqZsIylR
6o37xArJRrY3xpRYh6BUj8WwCkrRNvT3wsQoqf8Z5XKGSvvR6duAJXnW+/7YBPx8FzNZYru+BnXw
ruuZD/bzYwLR9NBr5LK8Qgx1n54NPWosheFK49TEA5WyHt4A4q6WA4GGVLqu+ZwdU3W5SfPQSE8S
voir0LOnxppgghOgk9ZsFL2gbOtD1fmJFTQ6SV2EFVZIzqpCzAul1EWW1DQU+7Pj5ZeTXn9MEg/l
ZYeCMP1grZ698tyseV4AenjJa/8xxFUDX83CwhVBnsYSBZx1X98/O3Kc6yLDCy2VMIgFYF4GoS0C
mAjPERoxoe8QhwRn8xDIcgVsuPdyNwN8yVUk0EoJP8aOZ13r+bMD160RP6TnpprpygGAq1R7EgUj
/K4FdO/9Oau719oll4NCdNCE3TmiaiqdVCKmWsItQ47cIBKCDFbILj3jRx/mYaYp5dW2/Gyee04O
6lHZIneyeLMe7sx9MHd4KsBjpZtmWjyVsn6OHP/QBZJE2LrsVJu+hh39gE5ibjod9MJyRb7R4CFI
4V0hLkzJWMohhs56liiwr2DLagTXxPJDEgrFRnbJsQtu6vI/c984IUPLDvQhGCpZwHS9ngq00Hb+
HPOpbhbejag6qC/gJO/H5kv7K+K3a14KbBnoveEJ7b0xAw+WCvgM1FdB9ZeKSTEf9L4LsfdBiHV5
DkKOz8YOHx23tPbVog81Ku9fpLdAu7FBum6jNRkfYh05hx2SGKYc+bPFFj8+Vyy7X6FI2zpUmuZk
iky0EkmsmsBl9kUSWxaNSZetV7JIRA8NtPr7ApROSUC7Mv62t42CBVxXsB10Wvs1UEdlK83BxIu3
4922B0H9is+PnubkN2EMUtY3GfmFQV7+pllS9+Tvm5BLcrkuOt1z0zI3hZDaTXNDY8hrcqJ26NXF
8LFj8m1Iddxsb8Cj8lJtNgrl2v0dG7rdg+VgWAxxCPvLJmtRNMu6MFMSEHpc6xZZ0EQEV3WTG/nt
e3iio2AXKUiHVgyGcF3AfxG7Lkklxi5byJVodYe+hGttbbWOtgJGnJ2HYMAARe+73DnTM/shyZYL
hdDehO42SUJxJCGeGTZohRvrB5EBOe6UHxyNSIwHp3WMeU9vzPtAiaZBOasqE9tVT1lRcMt8uH08
QOGKhjDkbNI0Eih11kaF26b0HqF2dr51VL8gQ82eb0N0NMc0x7+XVaaio4pQJFVz7LOLVDCUMbDa
t3K0KK6sBFJwVkH2ShB0mAhF9F15r3HGBk2mJQlrHMo76cOloBH/ilaYAlaTkRFsLRhBjeGIU8af
eeAj7wighQ46NTb/95mz5tqT8UxcMvvrXBrDLw1/4rCMFGBGIM4OlK5mOoEbp1eDg1gYwDGHteoN
QxFjY4Tr++WBh49+35rsxhVNndpI0Ib7eRR6sUuKXKnYglmlqltleRTvjfgGA5UjpbO3zP20Hns1
/cFA7XISRLVvuwNipAm2MBYiCNT6g+7rGcSokU82B3K4/u25d6flIlEc9tBVm3EcND0Y7luFlExV
/l5ncCDblmk16XgmaVNZM4vg9JeOUZjHZfX3znG18U4sQMSse6UrAyPJrCwQLa6jgdNN7Xj8yddJ
xqOkpDt/LXJl6QOrIY0Yem2ljh0U4w6YLEpKe0svDJx348PFh9jgN3Q7m5vhCMevI6uMkcg/q+OR
u54QavH6+u8R1FaSTvLj/TPaY/dyY8Il95/eBXw+8yaaxtH4K7JOsvbj+o4ID3FOoIynJlHym9VL
F5s5E+EzhrbiDJix+GbF3/RTBguy7nfGQwA4+Nh72/ydALA6pjSqxa6h4ehZ9X9+cQBoeDzuek8R
MuF5SY9FhCi8E86FI32XWQwFE3fbuJAyspSrrbGuLqZnwiMy1d7UATC3BhKFiLp9wbiSo7TCXtHo
HiiyWrPpiznZeeDSdD8OqmEYqbJBAPHDYSVKAzg+fbuYaRe+K0V1J7fRLPBqXvsWChl0um+kH4X7
c+o/Ta0h93Q+pVEG7SN9N4EpHF5BOTT9tgVf4AicuI+Y17dO//cvZpkp9kJkBdi1Tk4u1ncheVNA
yWE9u/SBj9rA5FXPBX48CkOtwOykFOVQ3/vl4369mbH0VrUhVqhhfFk/bDrxiZt+gBqQBXkFh23M
bUkTO+ZVHSnJzkKGkpuRna7vx7Zem24FnfM82APCatpruKGxBH+yEIkGt4bH9LRDUHAV1izHfC2a
efIkFthmZjwlWDqtoJr92Q2Xn24p+wzZ0+sUs7KwOcMSgMRmhGw3XdpfNSQg7db3nk7hIW5MZkyT
lMUZfco3zeultX6d3NVf+78/Tglk0+DNX+n3Arl1KQLoTuMZjs/IQSsDiNoP2iAmw+vwFpXZnE7/
B/s+Q3IeWf2s49jquFKjTDhJAtcGFyc0dCIfUFV1axNpbsrY3unz94WN9XblNltjcmxfqBYqmc01
nYH99b4NXHD4ho+P//xGaqK2I1/0+naBDGfv0IZAkI7kcNfAJgal+OvURPDUYlMcO2qZ/hZkJWrR
/zXIE89LaKv5NWD7bagtfVRvZrhMJ99Jt9zfQ5NSTF88uqcJx8ylITAeGxLPvUc9XokcYlWhSq8U
1VnirMHaV9DgbKGhw2ybwq38YhrUrLJXNoIndycHw4MzQSJDeNhRfCaFyBvIyQW7IePHKdpXmMi1
ytmX2lyhXlatkSUjbwIXdUhw/CzfguZyQtTENQU9hWTFgCWvgeQwRHllkpNrzU83mhUJBBq3ImIi
0WiihVMpTv//3ke748MjLi/gPtErX+QhSlpUBd72BZU1yatD2dPdpOpyXhqweNHO/Lo2b74NC1AF
dFVFOAW6MfDnbmWQ7fL5e7eSvRe11TEvj8j7T+QzfEJSs0TQlR4GoMueN8zWKqzEsNb8gqf7DQOF
GOe23ppinRXpuktDuSOezTjTwazt8NWy9b7rdgBM2NaFN4Q7yR0wleYX8X2uFIW1Sl7a+QuWIrgj
so4469T5V5KiV0FBu5/0wEspIFHIuYn7QDbdfyTl0bUU2rNVINTeyY+y369OgRPP9eRDqUnx8F+R
JT7Z0DvQCOAuSQb6eGIDo2ats2n0BhbCtSDIjmSqlXnL+VkdiqkyPcyUkqKQyAq877L4g+uHd49L
sSwU7lYZPdZfdfpUIveALN0uVdP5O9l8UNhEjncXZizMuUOy4pbwmUESJkO2nKEkDut5/QiGT0ud
+UfRMxnNEjlERQbi+cXjt3JSUHB+x+v3a+q2QvVUCieQQwA6f6JAyhoAiNHCch/uzHe1k0l65Jxe
JZ8R5tvGE0kYGB/gxDMrRLE8ZG+8Emm0df2c8cyp81GgRiXm/m5n2JFfnXsfvsK3/lYuSA0NB/73
URj2eNjYxkRmip9OpKU4IaBGoNbSdquujfiz6vZ84HkzYo++WODJngNgnvbnuYjt+I96yos7bsZd
5gj1A3zwRMyXRc6Fxa+PGth/r/j2O7fk7PUTm0hN97t731Soe2PMXzU4axbBZUlxHLD3rqlrN4NI
hl083Rh+QHcU4irMGuFM9LvX/vMv6uxc2QARsTyCp6894ckI5XHyALqwbdxq4tuDdAdwqQEdOplZ
XgJoiq1mN14vdlYJmgnns1mT1HgLxImsDgTDct/o9AqoyHRzD1UwQRd7mXS8+L9YEy6OXOsoFhi/
a94eUrUtijxBAqN/8qx0nh/7z0Te0WCnJc/sTULWIVHek6XhEshBFNjTgxzNkASBUAsYScF1HcmU
RPJzSE2bj/C5kWimx4BcE8hxVP6+FqVKxiaaWRM1IjFHQsQA+HpSXyRaEzKClS3NYblTQnkYoJjp
iUMyN6seFpiJmT/TnAa/sKO+CIHBM0mNdPI1JZ3yS+xagVBEG8fNm643G64zXNCSB1RUYawg8d2Q
EBt/OIjNcjJ9clHblUwZ+Ll6gYZjsbcbwcAejFhNS2zqBgn03oi6RxcjnXKXg6DZ3xWv7FbLrNGL
ytstLrC6HteowALyzxreYirwygu6wXnD9wLCxBHUmWG+v6phbaV3KlAeaF0OaiyzKfDVzjaG6QD1
DxJlOX29YA4V/Oa+Op4uBq6MOBt7CgV+rGPMLnjrU3nEI3COd2hh1nvE053EPhbpqEWr1oPAvjI1
QqhrijwJz4rzmF9xBSj7GzW3Ex8yLYGaC0ylKUqN7AYHuQH+SNkLfNi55Dvt+bbAzDBFM0jAGwY/
y52WCzWQh46JifTZYpGA6kZXJ9NKc27iA0keptUqANUOFImonWR8r5ftJkb3lxxyvGQOqyp5PbWu
vNdZ5CPVQFxXIMZU6f0ykIlCySScc+1ISkE0RODcKTft3DEgV0DiEgHQd5JE6W5+xHOLAP1TrDfk
hv5klQ54bZUQuKjIKt4UaZjpC/lhnKrd6/2IwZkQkOmmKtJipPcIe7VXJBO6D+6OBUpa9o7gu2xz
JQIjp3io4wtz3IZJf1Tu1LNwg8r4tDZgcZLBnWYY/LZu9IHFhXQ6v0fs/t/qrvj/UYoZedPIoPS9
ugmm/3ZJEWDmHtl9zae5L9Eb5ii2LZLz5juoKoZoZbITWvjsn4wNpzX7c1oMVlkNuCRmy7bqOexj
Hu1Tcx60tLvLh6Unw7svGTD7uXrX7+rWXr6Bq8U8CiYJeG3jPrCI9RUQmDCUPt4/Nu6AqCIi4C/d
AwMaqtrHgOxVj7d1s6zgqFVRmRS6c/DGFUldUbYk7gGQsnksWdzk9BESkem0+e4g8w5CtlOmLsev
P7VXBdLwUq8F7P2y1Ap/FfhkEzfKOleon6SjxjVnBVMk6NFSLoQZAqXaoQDfD22B3wjLHThVD+sC
MCs6KNcDl4LCLA0hF75Vb3DLdjpIyQf079/Ydf+SPqNL6CPCQLrAt90IFGRYMc8s2rCdPp+rAmOC
kKxNvEXp0dZ6ifFLyAWnq9osL/Zyvz6SjpL+68NyzcE5ABcp04q2SFUHxFFi7tQRqvXu4wyrqIVL
C+5rfJclDbJN9lFOTSGqZWykdjszTBk+uJEQ5daqQ4iUYua/fuy0QaVaaKxwFLfCKuz6J7rb7mC/
Pepp1TtmBtabXFEHw86Hbl+yZntk0I122i3rtLzvQWYh/5e3lKYM0wJNSw4nATUHMfOx6amzN8+N
S/SFk0AGK0h2nz/B5bQCQuvRNnt8WYQ48dJMW06ERNoT+2l1gakpAsFfojncDIBlc2oC3lPGpyg8
LZqQMCdRqwkNVOHMCzDKYHx71M6Fdf+MwwoDNd0CEhkRU7E2Vs7e4H6pmBReNBDBp9ApDmJw4fFH
aMWiq4+1zm4JujaC0iL20pqtzpoQs/IIa/htb1Zp6uP0WbkuCZm08M8d9HOYa1xY7oMbnv/b83PW
wsCHbNebB3O9wxsAOoecd0L+x1+FcAzrIJLJ6wEQVlVHqB9Wt3Km0uq2S1NSSBAIVamuD5mqvRk6
mJVI5clJg4OFMlajArdvcun7Go25Oc1IlmtT5gxxAgBhCsLKXN/rPJVTEBBQMqXSFVTCu/ClQ3+D
qDESTIij2cqlQaPEoew1uiSh4QJdFdvNLCLGUlVdiusKarX8z5T0SE/2MOFtre/81CwQ3XobXlhM
bOJfLRibjTXBjXFKzcDiEG/Az8FV3cBl83a+DVt+I+6SnxKVOgZz0Slpe3akmeOCsgQg8NyyWLnm
JsKlGjCWxeGEwcWao8eEDn84phBq0NQgfE75SQAwSW1qTDWS5Kz7tPhxSn8tcjCPM0smkk12XG1Q
ZMnwsSsHqCA41eC4nKu2htQVQVwNzrYxvp4M+44rn/UPmnOY9LqBx6kKAM7miRmpHKOGi6ZmJiXn
hfMByzgR9wrd2+LKOvmOBbyslTaCqbasTh6tAPDs/KIKeZu7AmxZPOwF14F+BHVi77EO7VPEoy48
ZCTs99Q/jtzGuc7Sxce+psPV0Gge0j6JUPow2Q5eqaMfVrokvAgfaWToilSgc9bjqpIrebOqQ1Sz
0r/0+5/BtP3RtBqDDW5Tfg7s6DkVlVPZ1XAf4L4RGzXPagbRnhV3EbMCnbPsdfqtvbJLD1A2dq5M
U43MuOLozARzJMIQpSIugaZv/4/wLCpVAUDHRCDj1MIjManmm8+QI1V4YiX4CscAJVDBbluKYtWg
cSkMJVmWI1S70t9ykIrEroVv/Z/0GiBFG/z/pnFNnLRSBcNGwV6C/yuLRWwBtrpBgwRjzxPtuebo
TTU8cmQks7bfx4bDhznUMa+/tPJmZrVZXRM6EzaxWUs1dxXOIMvWsUkDkWDvPjXPGSxrcw+iSt64
WWeqLXnuXqAbF0EjNsIdSaZHwOumBBTtFOhKF3BNssaUSUiz87N9tsYrw4hQtVvPQ4HXdJurys8H
fxFJmPHB27OlGkBOc9rGqqpaSbKHyT+96gVXmrmegSlvQaDYWDGjwWxC8whGTkXYXuphzTGfN5oG
ZRietwB/p3tR62Tvj+R6mWxxsuGbyZNXED0yVrrAEACg5X/LDycEaW1IE/swh3vJDuIu1kBL+7l6
ylqBSWurnkOROZ2tYiTVrEUI+bv3KpQZ3KL3jEffkz2OC2v/tItWs81jStc3eKz2umKvwmfkIQz+
gEZThnqZ9IJJBy5awbPBZ7mIcyAQwMK2ZgLz+HgohfURDfwXXL7x6kSubDdhXaHCqRoSAf1+uSuv
qVpNOKlQ7138iIKqDlsKz83cdJD0mqMC2M5dvDJ4l7d9JnZT39EVYHlLSnVbIK5xpDEcL+T8cbeV
slvbhJui/GRWUMT3g2j5aP90zMA1Wf8DZ2N2jk0tBEQ425DuFDhQWbc3hXCCnxotYdaI5IycDwhq
cZV3BfDT2XBk8pA+sV15kQ/ojLCR6PLp1LKjNhLAuJWstQjvoRUAsDP40YBVS5fjkBNlD9yT3l+h
M7un0hah1dXxEP3TukJtCC2c0iT2HhqOeFltNjzGWJSUCxk4h5BY52vmWymPWDtPNPjnAQpJU0em
03VOYAFecOhVQI01nxH6tbX+iqZb4rFTl0wnd7A+oi7DVvqFncuS7ngIRZTnQlQL5gskqda3GxPE
P0Ne4v78sf5n5fttNbL8s0Bmhv2W4NlGkpUdZf+Ck5zF598lsPYuwE+WAqCu4W98TU1yM7xv3sFE
L++vFSTgmK1QtN46NjkR9AmZ6/yHAtA/tibLbH1hCgEN/405Ycy8MZP/c0ZIdVNbyzVwsUwku5cN
LFq+1XZjq3/7DU+fkPLMUZG4agiNRhB901IS0XZCyBr2VZZx0hufVc7Z5hcUzqhCbGbTLv42a0GA
UMdFEGOedbfcMJFMb/XTHO6A+QBGkJB18DBcLrCrmjgiTSG10IibsfEizlkkqq3FdUCx2Pcg/wGf
X2dgIqN6bdd7pE4xyGuukb7iNK3024339irUq1dAQQsQULUqVoaJO6Y66jlf1t/lpl8iDyfYmuGH
BbpLlLV97AJroaA7eRWKt1NDNvb0J2noGyoQ36z3Zcr95u2R6kgb1TMI5+KePeWuSYFBHJX9QkbG
A1k5tdQXV/JH8fjK86KhcZLMMc/lrdzdjUVVfWpATJazI9S6/UeO5VM1efS+Fhdkax6EcsC18Rqm
wIsnu5HeWjILUHO1Rnn5ENXVcNhu14b1iwTcn6VBxhWFAnFcaBHlfv3t6WKOtk7q54uU4NhvA6/z
LR3Dz1My/vHr+gQwIoNrvqmqHZHpPzN1fqIb6wu1vKshS6lqfwCpT2+c7uxyio4N5xHC0xphu9x9
q4WhDdC2OBgRelUL5e3vxJ6VQ00IuKZvE3zq0Z4U4cWgkjqIz0UUnJ/ieMFJzhQmHdwsV22nZxpC
FYQ6ILlN+0IrDipal6sPHnqRiuVBv5lZ7NWEVkSKiDHSoWKXAV+G4nUGynP9VI0vZGjrqLHcuQWX
fGwdz0eHR3T55VT0rRZuXcT59SjP1AgKn5zCSZ33dpdxiA4uOnMbhKkP0682Vm8TOeFXKTzSzlFy
LRX3MiRTz1NMKzSpVu7/OZQ4iosxBLxHGiHv6qSBK2fi+nEjaUZr+TPKunKH2be/T7Jg9ojs1HAv
jLIkMgJdqPtzmNMUBB/0tF/rLuGgCda/DAG8spiMVvnrpU6xV3aKQhJc7BVmUR9s7rqM4WLzjVy2
bKGG7dLbM8i1eolnWBEACYvytKcZEdb5Yh1yc2BuWlAhfvkmXihn+uJX3xoWT2DgAdbt5zuRASPO
mYLiv0+CIIFA6f+ApNuZj+oAYjSFyEWv/xSUEFYyy0/6gQ5n/QFgINM6/7cJWKEQE0MbkNB0xN26
xzPdp2njhjugUMURpu8CfVwGri+6bUd3OSWDD71qk6qtAb2U0xnnFNF6mCf8a7FWCNMx/fLaEY77
u82Njk3BDDHSWkyMukv+Km6cmtZp1/HiA/MY001xwhO3+0ZcHQGQABH+CKnrqZGO3sVmOwrExTEy
wmII7ffwVIIx0XltckroeHJhqDpaydLv/p3siHtqQJhYC+Izi8WAZII3gzSjP2mF32PtEVbUae9d
OZZ4rSG+ueVNYEH/czDT/KLM+yty6AVDoNd2L0gFMA1lJO0MpkpIIQks2Ce3nECUrePN+7rlYsqQ
HKj3XFDjsnI3qExYAoIIKYpmPuf31c4Ibjetwz//GpROadx465Uzi8I3vV01ksi934bA3blE9CTo
5w+IiqsV7Ff7jv0D2yDeellk85SZUIgV3iLk9i/OluIQhorU99vDcf7w5BzS98/yRE3hGItQdy/5
7kyyBMXDlwF5s0JMdyplwRTnw82AlFCjyvAr54BLxSq0D3YyrRaGtqOmRRwQsEyposlDFv8qYzZ3
GXu5GpLKf7BwxFDFuFjiMBv97k1oQ846V9Clx7sflh0S6Syi4riTyp36mFVtN18OP62/N2WTajn7
XH5ovbuz1b35931NFTIDnXkxcMGw8DAtuoUoGSPRezofjxnXAHJQmGWb1sYsRW7eDZNAfdgFLDQo
pB/rLz6DIJ+oxgLahRxflsrZEIAcd3tk+Q5JpYsUruxZ4G7v/0UWKIZw3EM1Sq+oR9udxKQr/7wI
Xzg3oeVz+Wo1ODaL7ojRJHGKHwVCprvvBfkr2V/VPnDyZEFuKX5nF+5iNS2t0MGHSLud4qEiUccd
cQKFQ66uHaXLexh+PKSC6lc3Ncx+s/VAJmsBDyF9dSNno4YkaVSZJ+dpniyoX266lxLEAanKX0od
iVIg9yLjyrzkxMpguvFdY+ztLIdaJz2KOjpj1wcqI21GlpVQSYJXUfklSNUnO4Z13hQLtPkaURQb
4+jPTA8dUhD/Sda9wVxB/pIKOCsDxolzLHhImjXAqbcHbUAOrsbmGHvqZgOMqpEF/mAaWPWPBfL7
ZxRCsy7c7cvJn2+3Ww6Ceg9sS+mhYgZPyQnWLt33+VpJJf6Cqo2LXRbiZikkzGrgoeRRBDzjUqR2
99CnAMWdmNXj+iTYa8gE3KOhZZHTTkE4g/RvhEMoUCy5PV6t40Bgg3JQWo3eoxImXRY2m63Xk/mm
WYMS7PpeaTFczC4A6XhVhp6xcCNXrPTq3ptUl0enqtMm1sX/xHcKjJPDNXNOtGRVqgvTTjRAPQiZ
hOJKwvGvbd4zGtSMNjT2YVLzGgaMUCFVDZAeVa6Q2I2MF+BdfsGPEdbOMosFp8VmeEX+9VC9FNwo
YIaZlOXbE1E3PYt60n9Bwz8f+Uqii3jV6HEE0cIdcviIivQTGLO7a6/4Bz2ii6xXoOFLdyLD3JmG
ePjMBV0mwgM5SwQmboomMXD6T7+QgckxlY29FdwnP+URtkVnlvne9XPQ39e2Bz1f0otLMfiAfDbr
h2rSZRYbWQupD69Ue7iLr5k3J/1GrfnBypJU2aatvecHKn7jAOW2WlG2BcDxrkcu88E8WcHi3xxc
IFhUdo5DU996jTbZomNZOXCnP2IfNwyY/QtyZQUXAjpuFp0bv8Mnl01E4OG24PNQhPuzJ6ui/xBU
Q08pgJh+TF1s8FNg7nCEm4BY72helIMywjZlbpd/mqWXPJycEqD/irS7uQS7n/k6Jre2GTpcj21n
TEJ36IJCUnYR6wnVwz1SPS+ld4B2sq+gScUkLnMZgFWRiZm9yxR3xlsvrZ1lHGsm+ZtZPxUYztma
EBTvDMHLBfc4bS+6+TwWO2qxDzJyd2F9DgiIePIMMmJ40tJM4NqAzaXgzNycDjXIa+4QSa0EKPOu
0K/IomBg8flTSEGTPNf+U4aBCuPT7rayHdtpt1MeTzyWAc1d17HCwUEdS/1SPnMmzAohxEhVsg+w
UiBffQYoK4CxI7fsAPTeRlPCPJmf+bYjq90INLXvxeYPVhgoSgYrxHz9AAAHgmgf5TYQ4QpwRDB0
PVgk6t6M1bE4YjYCto/0xPHb2rbMN/29Z7JfMP/bpimnn0EeR1Ce7d+SYN725CfWQSHDo63ic5wD
WD6LPdIYXXMQypZ08n6H/7JkvqTV2LKUdkIJ5CChhaEVRRIbSP1aI0XhGIDS/Aan7i9PiaQMx/Bf
STIfQrCduKOdpfp6WfaMollzyz86FHzCaxdoayQdCtF4dat6t3huxrv9U+T3e7bxnJ8gM6z/mPy8
41NS0AkNJ7Hc4zhftleaDa14atewdh9tf5ND/hG86Ecpx9Rj2zatVEzAxujZP/EmH0uHy3JtOQ/C
cdR4qLMG72kDZmoArI+idxdceqOe7kF0lQx6UFhxugzbRYIaGaXnRN6RxjtQloMPbDQxO/ihOXII
K6lW4hMoFnEi+EidRYQ3a9tyDnT0tABznU6NsxSgZ12s0KykeTp96lRFCqn+gtv7z73wavU9w3L4
wJwsErSTX8GF+G0NbJR3C7vod+VOVxhlJqnndR7fmiXHHUnIO6rU9PrRNYqzWtjhimVr9ZOBUUmb
BjZVTN5X4FyyNRjLlVDhlgp1kcmZTbrSRBy+csVR7gnmO8aMfD0TAnOgZZPViiNoLaJKKBDqm+lr
taZSpsnVRyVfNJBC1JGz2did04T5tUca5jvUJTsKTNlg6MC6IfonV8lFklg8cW/Hth1eHNO3OgQQ
il+4HSAZi+ToO054opWcD8ODGuAR7mK0JvEOlArR7eNMGHVT9hX6ORL96ZqhCAn5UN/6K51f21+N
5/mS2jiuJpDhatW8JkGL01qjMLP1AB6b7Uxh5G+fAKFibrZy4dziQO861EiphtZJYkbgIK7xOTqP
T7ZbtqceJkntPNKDIee1dACOkZpHjUgVqhHp8BVGd2NmwPkM8BV2txe1Ilk3A3yFyA24xHQGxa/J
5Ry8znCQ4iTEofdV2xJkJ57F20LGRqpWg8PnVbUAiJmKH5k41rFBnl4KkpX2VivxLQJq1c1dpmpB
9UV/L10Ax6gBGIkEdso5GYA/9Ya5JeNKoHvWTmLylIM1PqnaRoqI53omlqjajZ5BGuZtHn/vIQiy
jHV+l9Z5eKHRkY2cpuR8a7/R0ulmNLh6u6brwo/jp8jyethQLVbdhoStW8KG0n0s7itnQuVXOo/F
qQgfcJYMJXEGRkLOSPgI5lY+KTCIesMK9lW7YDKF9aUoFeiWe1LiTo28HHF4k0+txfZGMWrYQx7S
qWDJc6kXtauQTP4icCRI5upT7OlvQNJJaTA/HVFG5Hdvd/ZXhGvJZfTvK/gll6a9CHcq6dXjv2UG
/ux2K4ePt4Ie7wgi72fl0yghFw5oGvsMZHdicpWsSQNTkehTTEDpY9gZ24L1MSxC5F4JsKN5c+92
7MTVuwIdQ0vV8Cdv19H+72rQKQgx6xsU50ddZ8qv2eui6suTHjHiycl1Dagu0HOHcDk9UWwggMgx
RVwCrs2PWYFUZahQ2/LNOZsYPYNaH3M9prWnQimUu78Ww3pcfZKIWTEGVaBfrqIV5x8VZfiOrSIF
7CMgKup5QGArg0K2TAs5cl9IY4G7TVV5mjZqXs8JZrW/3Uie3dquP07qHqeXE5DHCjQhSHhPB9ee
wBjZ7jyljFBAPgMVlbgthiHo7rBjyC3mUxucx+q0yKhBiwQYakyv6wjOGE462DMMJ1kDA5riV2Nv
+NzmRjk6UFLpqDf5Xy+1BvzuYWZA1zsmRpl+NjSdVx40xfQvJ41Cw67DCpvharaGbaMWGme2SmTn
mjbIhVdvjDRrLRj/NBc4vScgsWQr1JyaOgmv7IE++IdST1vdBv51cKnIe5ibae00rEdJf4fv24FT
S+nSUn1PWeP//Cx+rDSaZR97LtRRla6sI1/pK6/45iAXlgICasK4Y3oyTajdYG8E5LJhIpCMbcnV
i5Wm/LfUo1LoyYqjUTWdYWFeNWxsDle+J3Tdjk6zTN58qy1rPby5qAytK3EM2GnxYUCKV9si92d1
EU37pC4rr6x3LG+bWfRQRoCsqg+OqIIoMKf4LxnXEnO1YNCuIvATAJvoLbsOQ5ZzMX0vLPJL6195
XKheZ/akuHmJcSYTU54bulO4WUv9cm0LyfKRIgfJsTo1xngtwsGK1IA9IUQ9IJMWAXfQ5RKvgL/E
gkl5S4up0hbyGXh3NYZEklC9eAXAIQ/fUipUV7WxPMvQbQq1Mj9+SrFu40/AXup3Rog/X2zzY9La
g9fBHMPyLLE5E+xSD/oS2S7/bnMkKronQrm55dzPsdYl95oA/pVsQk35O7VcvWspVkp+WUwjvdpd
cxkiYFLT7IxUnE0sGgd1+gza7sd6HEq5SD9ENCxeItulgs4tUa/McEWFcY5q2uqcNqOCjGOOnHyp
ljaUFtSo5ZlPaLJbsRCtEv0bjYuC7lww9tZoPRRNBJCBxm+P8zgwArqQXrlamsgK1IWoXx1pynZy
ttDFc7HgmzJpFc+P2P94iUWz5K1EmOi/mefcu1mrrFob0x2ZwhwmMNzGLRu0RvWWgqkVUwjLzS8K
hfwvdXi6kdbrUiztnjkcH6F4T0O8usDLqXQQsjoSdno+hWo07zfg0saH4dxVO8MUBG5UPM/fbFep
Z52kl70B1LfkXnKJNXrMhnIiXW5zQLoncnvU3HdDq8ho1xS61AUoWiz+Dv9Pi42FvMRxZcmwRFOP
8r96vmYr79oFXDbBU9yz964Wk2HKZojlatDM0gICL0+hjI+PHKqCwPRJcStaqOdIAHPBS+Lm81mK
nxenAeBvAGoKQpm5vxN3EMvORGilZZPdMPtn8QB9CDDODMb62/UEc+FGYmxPC3pw4y92sTdNwmOY
4zl4RQf+JJiT+LkVVSeGy2yKtgDu4W+t9wS04e78Ey0Za0bpceH5ONnoJkT8hyAK8y3F7OGiZZHf
Th53Lk/JgUGrjkqxXv1DkXTGraShmj8pxnofT4ls95P59C+ujT+0YEEmYwstcNTzVHDp5AYxHSKt
gWrgdEicS16jKBnBlwhEFD52Fgswj9IXDBp/pCQnS8byPdV9Bj4w+29L0ihtF2eEifQwn7zpfOEN
AINpr/ltC2oP5fHIpidgIHczDwdYG0akcwVYjb4T4DqbdclG5Whb4RCumeYX7sw6FKyCu6mVzEkU
9+bTM6VOfb0QAWgNKVJqHBl/DggEvYujOemNCrAhA4rfzYlLGrVLlCKD0hfMe85mqopbENq5JBqJ
G1rm59xuftVvPwX/X07txRz0MAlW+lkB+PHOJL/JudaJFQ4UXGXFK1RkoTBKlXnaASVyZU5YMNdh
yG6sRX7oRc7BCTHsRYmwFe7gRYO0dNNVGiSrKxrCDLMj5vMR6ZWPIxpdmVz5agoWt9u6l03CqmYd
xCwRMMVf8FTcBewZ2OgoS5xRqTeEETYE0RRYz4+01ROvdualTOR2c00F6OeqcyvWer+j+5qeeCGV
Fd6jIMF0p/GrfEzE0NdCjlySFkHCK4zFXXzCKHYv+rdgygxOxE50BJXIY2BDkQxQoxvoCFTzP3WQ
AWJxsE1apADWvCxQzYTV/KC0p6NmBFHXA742bDuV+UO7Itx8ZnfZMtFsTCuIUhV++DmHgqXFitkJ
pK2/oUygTBY3pgU6mQbxwlXg2Gm/aURXzLLrOXVkk1VVASpReUq15Fd1hSxOgJCVlnPKRSBKUnYe
mqn3/btzj0dWtLKcFSMKt/lHvjpvWxjBOx46DoPDgrCI71uTEUs7sQBIzE4njgMwbW/VYE3YlrM1
x/MOJ+k73PxBc2oLHx5pt478e1lmP+1y848X9i8FHCxLRfqY3Em0Z0p72f8Z5oDhqsT3miEb4Utt
HHqmBOJ/61mNuqmJ4nmlx5BQpZnahPURyeb/g5u9OTBATutE5zv82nzCCyGVIOzs5DeE8PcD5hcg
VYhJWkus2ysNnOHY9crrxoWljMM1qGzZ2IhAXyN947R61JU5Ns0X+2DFZDyygR6s1vMQ9qQWQc08
NfVX96bamoAhgaSTli4D1XywBEgrXfJg7mhWltvodlQ1SF0rPm1qpZKXvrxKtX7E85lIv4dEzb3o
gJIuX+C3HXVo9LYoxjT/ybGsAKD16XyPrfZx5SNTR0J6/kUD6MIReO8faWDs8Mc63zqfH88ASi2L
rGIrNdurv6BnXbpFcVm7zmTJ2OF4xWLZH3HSEBQz4EMgxYSQDP3ZA3fNPGWTA/vx7HcNzs4Rg7Sx
Pb717tuQmgtf2PcCm6Y9fxacIjAsTfRgoNPDEtJgY5y+7027g8akmLG36qKu/ieQ21tCct0ijYoE
5vHeCJyYX6/V4w7CAVCuj5YinTqQzedy42Uzij/TzmvB/h0gKsXWBQL3lJjhqaH8npPkY1q048BE
UaQuxqgbXf1pQUA+27rg9E/5xfk/CH40VRIE/usifw2kXVGON1I4OdskwhfrsJZWq9c2hh6l+Z5b
agSWG40/WziXxrkjQGJcqPpUZP2qegByjmHHMC/gvAC1d+fnMyNjFYi07g4sYZtEgAaOMnfw8vp2
D4OT6Tqa9cQfMC93jKcPpF6T5wBJ749GL6hHiHvKCfGnUxNpJNokki2ngoTWjetOCtc+fyyH4MDn
jUxgXKIxYdloEmtSNrzSESiGjBnq8t2VrMXK24dfOLdDglef8um1tfZBIqLaab5Y0AmseIxxMobL
bHO+if2z/Vagsmt9+JfmoUOKokzWyxw+YH5dZORlMCN9y0U9LtRO6ox1tcwAseeRtUpGqRrCw4b6
CQ6yTtOcyHQ0xm2+U+zvgoH8HEt1MrZAAyq7+r8PlsOTSEiv2CQ3h4/8poodfe1Y2eP8xFd6wL9R
MQtP+xIx2up8KgOOQM4OOh/pfUOH9jexWgVQpQX5t2bBqzuaRBj5ISwiCp+TEbl71di0/mfD7aIY
sQ0WcmjS8ZwMlxp9FXLlanQ9eOybC6T2+BCL3W+1Q7ArfyEfpBxCGKDuX5hCLIm/z5BaAWRTghXz
V9fqcDREpJA+QtEuHzEdwbx8y/1dCkw5yynoYqQn5b1IF4EhO6Ia7VVDxKE75GJnLI7fxNeAeHi/
aM+6uUuILOa7hnypLK1Os+2BIzbWhoRuuAOCfZ5dXpcj5TNOVzvTazsWOfEpI35Xa4CzRo1XuqEr
Jc6zzCYvXwBn0U+4YMUkWxCJapP4ClZP/kgxtTODIvaY0IQtcGNGD8n6PQkKQzJH8SLYVmvQH4yG
CHnAqiyND2EKNJWsBrl3ThsTtScujsHHhEvwv2atQ9QhBgP9oJyZNZUjs0Gehmav7J1IOJejNZw6
DcH9wLlcyTlDeJ55Dce9C2IrV96rxohXLYWwxr0EVYkkDSV8gCtpyPeK0pmZPoyrh9I+d6I66Pr0
abQjZVDaJ8Mq5xmLiRgnrH4BBRZmbVHT7yfyP3wFueKgF7h9fnVnKUTOrFpV6/Y3C74R+4MUPqt1
HkKkaB4t5g5jiAV3CPr2cWCON4cubYGNvF+wgPhRYPEndcGt1mCB0PUGMFKLEbRI8FCLhk8cF8//
Lu8MOTY4CWWBWluosIOZH7n3AiYp4Lomdumrw2rf3+jrIuftuxEcQDQMDMI+dKVWJo1qnTWQpxxy
fYLIOrKGgVkdGs3C4SwGaw6TQ0/28XX6E6hMcOnLNWDSc33gM98M/Frx3wJ1YMiWQi3YAxSi19F8
mqjAWHyD3ywiG1yyJAXWQZGHNv3zD2EFBEOHDMw1miFZue2Ng8+FL39fBIJ7d3JFYzw/bJU9Vvbo
rpY+QB+N72pG0Iet8jqWK5wEYBzJRjylT/yt/+EtO9rNZR1nbEbHYLZTFJStV0MurUi7+s2j5taJ
wQlTRmMmZNYVciJJQTj46zAVl9KxBbCwLLBWCoSVeCC9KFNNYpE/iLWI7DO1zrVlw8D3oSE5r30b
LkdeXn389r0IHY9p+OnOnar4RqnT5domVK5jBYvtHSJwlk4bhjis+qaCo3bxmwR1C+7+824GaXiC
e0uEkP+FMzbsQ7F+jMqQMpObCYKb6FZEhQJSrK1RZ6CTCfNfRDARu6246ovmCCjaZ0ufEBcl/SmN
5fpMTndlcZtXmQJyC1sf+fumE1BFYDG+wKzAjxKfQXoFvlMooGqSzzNex6D9r/89mt8XawsfM6kU
H+ozC5lharUyxmdKGVyPzJjCXeHMhNn0Ubv6EJVDRmD7RM17l/FJGx2W8M2J//VeMoexTDtV6jIJ
GAxudtCO7j/aZwtM/IZZpbJe1VOQHr3ClbTBn9fgMLndXtFqztoSn0aVUQHjYAu025457KfvANCf
1NmATFfwzHmh8t2R5CLmtM/pE9Jg+ksxJqbwlMyPRGi1GnxxKBpFHIhDmLO8C6R1hrK00bgo3Bnb
ze2+zg0/P7TPJQilSz0MGMbmPrIsoxFakAur8zy9C1XKBtmLbkTNGATl7jfIxeBLnDiQWLir2VCo
v5qDgBuOJZBYrYLkWAq2Fq6eoC63VwyZi1QAQLebMH4gGKpnldD7W9PRIfwlXVRWU5Mr2IxL14g6
B9uqiqsHvefMD4Essb8ZVsXmSr8zTk3p/sgnpmJjlrKpLbjKWp4c2ayE++LpSgsJm6e6lPcaoFrO
qXUPYxGFr6LTm/a6FXZSzmMvAfrOa8C8pZckTwogu8L8p0HUkb+wLA0lEP2OJr+2wslkNTkNIJsL
Y60fgcP/P+r1bybYb822wyIjehHzpzsqhTz0kb81+qO8eclp0xstUDvZH0xiWY0QIsDbk5GPRTZM
tqR059Vyh8L/36yxtN1lJPIGK/kuU40cjmUFe0Sk1tUKXqmgkO8aI9MUza+SAiAcUbSsgPSklpuA
RFbP+EpXHQhByqmhr9Vx5VwfjKe56v96gzGyDJlTSx2d+TEvmrX/T5+54du/IYhUtor+9en0yM4/
6QrcSbcaxfLKRBxLKjpb79CnaE2tBJyDFJFOVgsuuGbw2wGyJVvq2CGXRMhgpbO8YNO7+AOA5wL9
cK7LlPzeZs+KIdzFqKopTXfVy0FICsEcAMVbPqLUUNfX+Sl0MqC3iDuND/qgtRw/DCbVGNemsujd
FyEpIj0Vl1rK5CzPuvsuaXcW3McTdZlR/8/GvUMfTgjjpWkVjxJRCLVxz5WNpszyloDsnoBsAIbZ
M6TuYJaWeIyGLX64CFubLcSRjhxs1b2Mi1lXqGtaNDkQRMjGBZh3/VR5IYOqTOxW9jDO5OrNpA2u
ZjtNoPxrX4X1BDqOQeRhNKGY+Zm1A7jXX+BxvscyqDM6fhr/ac2VAd+O+mmAsyYtuDMQ8969mZcq
IhszqCSAao5wmiLAz5sabfgVQCXlu4Osh2oLJskjTeq+wVfUQ3QKZP1SR5WyrVFmXM04UrRJgB6D
WPwfF/Cia/pxomwQNEGdsUBqX1vJMu6aEJ9eOwUgG8+dphHS1apxjoigkrFrHuOV+jlusXh3GuSx
73iJCjAYY7CIGTIcwBtBqOxmgXe4ggT8U7puksWff3K7mJCxN2NSmrFqG4UVTR0/DLLWSdXwGb5l
nqZESfq7h6Zus6wr3v2VokF2SqtI4KH81ko9RxXT62IpotwFyBnpIjNhlD8xCXO/MqaRAkKg09+6
ezSjjxus9q09Y1HTPXUaRfODLwXdSzGRd90wQR9/5ba1CVXMzF+N1INNWDvf7ngu6q6e62xyvxjh
Z94mJcMjb/SxXDlrtSzEkEGg6tK2LdxwIt5id4D6BGTL4t0PFBO6RC5/RiGWbA15Qd2UbXND95v5
bAMWaBQ7lRPqlRD+NM6CSbuxyknd7Vje7jbZgas+I+Gu/B8rXs2hha3qLSxZ8/CFhhmyxsK517W1
AsO/osVi+5Y6EvWpH9XKS4HZn0L1rb4wF2jt+1rh8zr9B9W05kLWbi6ey66YixIIixmRojM+DBxg
q5oLApiAr3VG2xWQjyjMtu787pqWGNWfxPTRe1B/Sc5YRh0wAv2arcIJTccTDHFuKsWbeWdlyD43
A7VokpEJsS0TKzT+vF+KayyxhZPM9i5uE64dkPdsf6y06nfGpBr5W2eC2xWF/ce5SP0P8LVXvLwI
PEdANdUorPtqLbj09uO28oZ+BaZ73dZyzpxPtsRzfrfl7u1HwxVrq5b/ZDnaJbs7zfFJWHas79b8
Z5OCuPJ2rgK5uWHFd31sDoE/nfJI4Nb/cLxRp8YKazBVmDtAuiEUG0OsF+vB6mefvlfaU0nPCiRZ
sgN04CqWyuS22+WGycVOgbnePIjhBO+2LHiOwV+AiNxx+2bfcjg4xVBGwsxvKzvCmbdbySC0p/q1
Ud4rdwq5dNmJxaG4/ZK2cGz8hQYQOePSWE1jMjmQ3oaJbnoHOD3+5+UdpfZ4NFdCKdaV8ndvIJmx
0Ln3/DNxLSykKVpjoeawKw9IAQr5bi7SKrNwR42yr4YfG1hiAsAksNWDhfr/fMbTWbPUaYApzfWf
NECPUDcqtZRfZ2FjJTXItGHSAaFOQVRJgKErirF69OCCP+V8EBqcfxg2/P+O1G9BiTwUnfiXhCR9
1zepnKzlGcsHKWAbmxL62fEGfw6NIXeoWMzft5zePQA4Biaq9wXDBvpbzVfn/VhZlhTUlqzj4KLZ
Do3bUAstMJQjlbNu1cvjZzGY3C0fF+AOjjSZRCZQY3sA8XdSPoDQCuoT5LrodTuAKxVd5RFBa8pC
b5IsoZMLO7RukgTojrU9E9V1oadWdWyHIjFjoWMwsbrSf+ksaRo/iENWqp1DtgMg/oVo/btdrYYu
FrTe+eG7mslF/ZOT7nsdh+Bartvz2cWWYbNUI3pVpO39jPDE5k4dRn6jbIjvg7eWkmnN869aO72a
75PXK108tZaTr/+5NhAV6Mh1A4cvA2LijpViotMhZo6pTVpzwm2B5TfHxhTZKSb3SMy1FEv6XpYe
AA7OBrrRUAuwIoC3i/ngFIb1Eqdfd1S3efZ0sMLZqcI+tTW7VrriN0dWDIsJaiFUz5jalqOeXENV
MixRRlDyIpNdBO1Uq9206naRH6YHQ0a1SdauLXXH8SQBBAiVRZFPZXDAnTsxk/SFRbTKcjPaYGRt
CLLGjTFZ+hytgSpoJ8c9B/uuLbMYrRFKPi7UNbLGlY+g4PJXplLEsAH8hOAEl0DUzZ30NTWy0kot
M1RQXWXtGNNBQ/VPVbbq2S+lI4pP43KRAaRM5a4tOLS8bobX6AfbEw7aETbBk2fNBdR3ezIExqJj
lriah9pjq5ENBX/4T1qGlL91e+Gr6aNcZnPM1Oa/yMG3M1Z08JxpeG2qQapZ54e9yzBEkHCvvuB4
JTerPTUo/WRbfbIetW9o0dPLb/PfRJG4lzczae98Z0foO9MLSTMdYfTxrSXEnk1dxkuWI8E3u7pR
iwQc3AaLDIuPlkP7UZjQShl2Ds/R1VUOsgwLXtSq/TGAbyV4VmMqAttUKcqAHBbbuJ9MIsmA3OM+
xmfRhK6d5fLTHlFiQhxkWre/y5dK9nStvRxViGXGG0kDupBE70WWd4kGu5a093HYTua3PXjhBlWW
1a9Btykm1o8nZ/apFszhpCNzZjdx94hZLABBisKCScVeYMUao8r65NYTWcBDQI+2T7JBDwsZATeb
qKnduL8JlXgHCMsEjZygPgurwJ9JK+l+SesuZMb6BP5tfMIbxs0UwU+kQzcZlwHDfdwWswVHubz5
1f7aFYyr1y/xjmHEFaS5MkL9PoqX+N7x4muabNfWxjwM0xWBWAnIyMYtaNUmSotlNzoJzv62tX8T
NrEfxHVnR752q2om78O2+EGUrqoCrXUKnhasfdyX+kDBZOuTXi3BTNBQNsiyHh1LPbYTt/4BsPV2
i6knOMT0pfCr2/Bejp1LQ+19hhpz35CHzAkVMDVnZxx5ftkzHUaLJSzAUp4yfsOuLjqK1BigDwPK
c0Ksm8Bmli8a5UpDr6z2s3tvODynydC+j3MNeDUOEJ+yjHAFVRBBRJJT8zdkFBOzuPt8iLdD026f
d67E7DMMZpT1KRinIoGpMwIm1nIHeIkIniBt54a/pQ9KQVFbPagX+3CITksG5X1u+I3BqycSNjlb
Rsdli/B0RhXvbjzlbOOrs0FoU60RH//NqW73UMF+3FEHEVf9dloTyLWyyYltU57pFQWJyjCejYdq
20aXlwBJcvVHzydSaG3XN3ngYTwzNNprD1mxQobR+IKGMfGe0HNFuhzxZ1zEPabHgRHBsM9oyuf2
yXxum/2lLo7foELJLXFQsz3lBvGoD4sMf45raDF+4u3BP38eOcpQvXjhWXObMTOe4NUtBGmVN0is
Fnbxp7PaOi0kmiqawOay+OyZkmeeurn9tPMbO5O2P/b+aB8DqdoR17gvOUnGDvdoDZxJRx7VQBYZ
95PzXH4xNtUqoUGMKHO/h/+uqqgzdd4p88w+OVVzJzRApG+GBpuZTgCxXKsL5R1DF7pxGpSL6qC0
vdzsr8UqS8nyGDOG7Z0ewPT719C5IPYsD2rbfuNRU27tZvm4v4VfkQuCgFTp7EqDDPdoFRpiEhAJ
bpFx8XstzFdcz1TuQw0c02CzqL2gPwBElsyONacI9vq+7HuzTelxuPbRXtYRUb+HGfc2Jf0mdlFW
p/u0NQrQy1xZA6iGIDtq1YiJuUBQlSjTnThkc4UNhCuNlYh2MgyUQW/V9RaaUYMC1pZKi70izB31
o4oaHUT/qMV3hV1ERNxgsPTbJL6A0aGzjYJ09sFDllJafp5+gVNMVGEL/S3m+IlSiD0oFJR6YgO1
lCzGjsYz+ixF28gsvxMv/CGDQ4EsJKZyb4Ai1pseO7jFWfxusfS+kLEExYwQSvWgNlX9OhzLkbFG
7nQFAxRT0oNm3xU5UYP3qo9gIEgG/dHsQefkpyCsQIV86bK21VoI15moRHWl8L9WU2PDJRXHtCXH
pO2Rd97ZMlk+GJ8OM94gd8GjYqk68U+FHFG0tOgzUX1NOY6HLZpo4AQPcTHjL5uB3owiv1Fr4vzN
54OdfkdjZvIo5Ikb/9zXxmapSJvL9uY2pxPZSXNdo0E+3fkL9dtRr6Jwk4jg50fOfM9xRioMBxBp
Up22NQsMsXE7DPMVBfEQcuiQi6nYc2B1PrOEKsG3mUX5E9mcgB+mnrWTmMCgTX+R5suveDAQ53DG
9c6yEjPkyfzSYgUpj71HnkwEQCsouPIp7e8X4TV+8vyNsuifXuhWN3jGFAWnJmpcvgdtSImBSWWr
a37Vun94DWAyUIOG0A3td0Kgalh6TwB2QQsZasxRxeEoLxM8jhH5iymBQ/LtL811fS7VvBzntxro
PQErUJKqLUn1GfH+VXDAxfqeflmxBd56g8rjGpf6O+QFBLrBeVuG7t+b814XQw6jF36wucuIlPuU
iHnIoSboZ6Wv5mBUm38ndozPb1t1cDV83nwZoiB7T1Yq8ikK4Z8XdbIN8WRwhDEzFET7NQokc2zU
ZIXaA7KaDmQZbNnm3CKE5pr4FRP+iv/zx37AE7jzCLpM+Z+rfiHu/kad1xFWOiIE0zRkJC/DHYbx
znylFQa3AGOf3pxWh+JLCSNdkhxq1M2fS9xbU4qICFa9+UV2k7QTfPJZXKwS3g4u8tGla20te6DD
gbyiZ+52KlWoLuEY2UPf78mrTf5ObRrAvwSPHypJRYPf7zmkv2HR5YTGVLWjoAgkCGw/2/zpC/By
YPqRRv9sY+apMgu3R7j8GeA1JDMWap7gceDf21AdUCnRGFcXfMgmQLEP7qBh7UYh3823cKNYr98Y
Y+nVB94+EQv1PwDVMVECw9bZ15dBR/TqEYvWgHz9boOhvpWTd02/Et85bqFyX6uIRmQzPwLndLiO
cVjZJpNs3Pzy19g2damHZxLrTmUk4oaGzgoGszJ/4Eaw/gFI0EkE6CzPfhzwIrlNrOHbpoL9DIps
U7lZUYr8UMi6qbnwq1spmK/DfI8pD7kkDWnsdObTbuYmzPcWPEprk1D/h6D/mTOr6UXMMRd94la7
rrZwU1YHPRoJuDp25kxraDpNYsgjI7mNYnjiqII0aGwm+WohmR4Q3lQmSBShelxg8DKHWDiKbHfq
lbvSiM4sxQ4hZEU+JT2lkURvGs3ybRvSpUWRqEGOAmqKZcT/YHPlKR/Cl3lyXZy9dpyFKT11Ie53
0kPC3AaxmRtekmtsHLHqLszfJakZnSBNulePtrnC4pu2b1Bdozblyr30gEBqnHMPlABBAdylNuj3
IxvEkDpCqjFy2IL1kdRjocpPmnliGvnJ6zamySqqnKTc/NLXS/vSKSSrlLRSSEN6eypNOFH4JBQS
XxeG9pMKK6XthdUNh3z0W5YOU9C0h6bRDaYI4uQbRE1o/69vwi5vxyOp9oMXRTtvAmEGEgZrCfRh
pemEGDn/tQYAMp6xhJBdMyYmpCawQsx/4t0NysKGQHM6i5xdvqjboTBKmS+eCis8nZAzv/+AQ2An
8JRbKYz6b5LpSogTOqaD4DS4Y+efVtfYCA1/4GB9ESJrh7W4ORf6djiSrVFG6C6rus80BOaefOZh
qjJZYZq9qean7MOIdGI/4a8WsoFS768snj2soshTr+8LVa1YigcECmmyQke841DuOBuyBzwwJgYk
aJybHHS1Kjo9Cjq05k4bScck9TnOQi6MhPn3XElG0Jcae831zSFdQ5xR4RgkrjHM9wbIrowoI41t
COZ4EK4RYm+bjDcK0bZukbrWD41UwdPLv4tsA/pV2aFrbLkm1vWcJq+WQ5GYc6rHM4InJpS0iOFR
TwcVlzloyemtesyD99C2jm7d+Bo8RoypyC0kQhBoPqBF0GRPqpU/wVsBCpFi8VwRucln+QMbkZ2w
1/F+EYtgMjAsvzt3SjoYFT+Ccvta3nQd1AVhXRPhBRbnin+5p5RBUanFULQqCSWFB50hVG6XAoPp
A5svKogple/JdEgTszHCyoFNKNBIsMPybo6W2tbUuWzZ8rKESnb+1gnGfw5NdZLcddZlCEwhoMtB
Vn8vnV0Q/Dxaf6Hinxit5w3VWKa7C4l2puROSHmPbefyGsG0f/163Ktb/1U9gqdvInIikRgHgKXb
cQ4hK50C83qoLFpx8PhFpC5n8OT91+fBtc2gtVUkVfKAfvPSR06xwWkTVQmgTSL8JuROkpoyqSv0
TUipkML+eB+GO0qzfbOu9Sn2j/vK2NStALqUg5BnLEp15g8KVxjc37SGB2871YzEOnAm3wJx/TzD
H3EqeFyUlJ7i50tXwcxEejs9+y+iJ7DVsYXmSvciUyh3PRTVs1wf3yBdEGc5ps7tsuvUjNyqybR+
HOT4lAvjKgn1Z51D/yUQ/TMbupgqHLmb/wVJ/pU15lD3Gi3OTDlLbLP3t6bb6stv9gS/rE2eLb/X
strSTkQHN2IfBgs+FGGKhl2uixlyNlAjfH1HpdhXPr/SfOj3hlJ/gW6MbWZsrsZKspfgKiMDGttK
guxspM5x2Y0H18mCR2/GwjuiWCeAVKa9XtTOIj6hRitHUCm01EI3VkK7e1uFKAkhe19Jtc+qEepO
8tZYvDDmpZsZBBc5nKRcakewtQGTjZsT2x5NexK/kvoJF4wfm41y9Y7bCHpP/oXEeF6n5iXH3J22
FgthTX81h449mWrocxeDL61+dDXw7PUtEdz7rAHioim2HXXftuJ2IBoFq1iuDu3lCPllYKSrKVna
JwfO9Iq0G29tmaoqIeXxd8Ve4eOcbcpZLPorqVS0F4fPLJTzFO/ttFB4jSS7cwvIEOTUWw7/u3SD
pVrT1LFhCe+zlWU37obZ8vhjJz2I9vTn8wmnZDadTShk1l7O+OZ4vXpvTzeHlMZf0obAE70Nc07g
OObh8JDp/Ws+ZcDeVZoUlEEUtfNMtsfHWFOAjIwp3OEWyqWE/EYvIhWvSbaYwXQYPHi9IQOtJvTD
Orpei1qPztjbIkSzSazsItJyyZCYal3jdyShCqOxwTveItA1rcxcovNIZfSCmg4gtmvGJ3uo5n6j
ltGtaH/UpYFBhd54pqW9EU6FjCDV9pMP2kjSHPcseSil2FZQ8JUTqwg8BeXaHdUUb+8Q4B9BZeZj
hb+35AJOon8SXmiPDScuOd8P53pILqqmbIcuBhtkKMLyCOfjv/zxzzn2I4Gt9LeCoLJpRVv+uz8k
m5Fa/frletpb58pVFfUuL3Iz6Ar432aNlg4US+KXqE48Vcq6msx80C2f2mvK4Re0TQ2GjoWmTi+4
lCS7wGdRQsaNyUzz4CRmHz8ThB4oGiReNth20T6pOIYs93OxlXDgNyrPBYQmxmOeM5nCPyCgooLp
2ix6HRfPPrOih1L/Nw6Ogrxij5D6T6uJukAUk0vjyCyJKOgocCogYyKMmEyNKgxYlSEpYcA2ZGa1
dErljAwdESZbOXSweiyvRtBH/SmQkMZ235CKSbEHz1iZFpRG40/RjpMjTk6fvisJElRp8VtYtxAs
zrBQY/Vp5KUd/ipz+ZB9mXUFeYEilXWf5xRDYEOKnWpssojMT3EKk+m5yiO5MhAbf/DNICW6e0Rr
JXNH75LerSoLiticxvtnFLAw2E+Mn9mSXs+gG5v6xLms3ww/7YQikeYwLZQFFDf/yEXqA/9iL8m2
YcisO87sBNtXAg7H51UhToF7y35ypjlxHgsCyNfjCoJuOs8KLq+PblMVg6lmsA65Cc81K3NAQxtR
A5VW+8mgm/c90kxgVsqqmQcF80ijHYd5Zt1FyUnFwUFlfpimvq/2Y+tL4yrr9TxTxn1uNbPGLugK
hUhoLEeOW+T17SHen/bqNUhipPkjI8xqnnPkS7a3eNcOKFl0e203ZV1/5yCG6tefXDjpESNDjWI9
0eSOGouS0AGqT9142voRhvSJ29czSLFsYqLMumz84it6XnP/OFykWnpgcen1tCWuP0JoWjj+bs+c
lErYEi8Cra9dlnIZfWjI5NBKYCUcmq79sjL27UkoeeBnGUQJNTOA8IXEnNC5sRLuIGeqsYmMZj/r
94HdPaca23rW1BLv2L+9AIm9HzjyS2GNYKuNze9n91pWxogcPjDCgf55cmBTTMPm8bb+/rWYuivf
MHmNMs6V/AgthhFnbioOCM1N0U7k4AX83JQiXOQ9VsSJO80406/uXW5EEIQ9PWTyyT3h9WSce7KX
OetF6/fb25ajBpk/C8hJGkYMJfE/TtZAQmxRaj5rTsjyq9V0hTyAyBCixdWf5rR7A8A90gZKAxU9
MKryZ4DFhQTR3EBHzRo4qh1dqdGMAK6PycjmjBlEGQ5EFzHEbfasFv3rE+r0/iWBayP8k8grPiXp
2E7yvSKIW8gRAN3r63EjmV9WOjVM4rVXS1u/n0r57SK3b4ybgELoQG1vRkW4GQItnvNpGwSshtAH
PMXI7mOgd7uJjLAZE6qaSS6Udi9j00A/AveL1pPANAv1Aj3DPi0vDEBVhMO5j2tIDBIK2DYXiLNr
ishr7sVQyZfUiQ5nQSO6ZJoLQHLnaUzx+4qODd3pHxXnb1o2HUvs/6anQ7kUXNxq6sny+Z4UfBA+
g4WgwQiUXq63t6K0PahiYLFot+qaopmrAZ0yfmUnM+fvNlmOwwiSpb6mqvi3rx2+QqEruvgMbO/X
U7DC0+aL1x8d0Qy2/+o/EP8Ou6cY58NeGJYwkAal3AgdQCopF/FQgKNdcaaws12BtckXCqD3fPY8
HZSJpZirB3Cwd/yF92iWwgQVdo6MAaoPy3Sgz3xaTDbp74E5rIUW6YOpBqUw2604d+KrYEl8fOJa
QVN9GbAFuQEOcbxfGcwQAr+foLvNzgPxJ6XMY9koT4mnnZMn6ZSDUtOEQteHyiTUSuKAHSurctCj
WhAlq2bQOAj+tgmpD/P7foHYLuCMSzmX0ZbR9Kn9J1cHFB+/monW76GcRIxB5jFEC+ZDjGxFuH6a
HGa9mHGPpjMseHWUguIySBOOEBumMDilxXB9d78Yq67kz2ChfOkAko394wG47DuYiRpvyJxdsg+s
K+84bUcOHo4nz/XDFBlUM60mjF6afsd2h3RiaseA74uhAMnrrRTg/436s+ACMNVeDhP7387O005P
jHTUQqp7tRPGKm8VJBGrnlKrNEv3XrJzw6qL95hLVqQInXXhwLvrQDzXqQC0dALHIYihZfoC5+pX
bncQQ9AKQ6O0+n452zHeVR1wROKV/GjxeGjcN8gbw6MiX1trNgVMjf//2hfYyTijfzBfWlSRvNno
7jtL3X/z16WeTpeuW29uRWhzFzIaVzshqiU7owNXJblINh3vAdcS23IMNzLsLzsr50Kp4HgQTNwI
BGd/F2CAiFVgKz4bEruCStMAx8cmHPHX9OuMB6x/YEvpKkZ0rYaIBy1klI909FN19RKhXBstnw8T
ioyHd7WMQtX8KuFJyhfZI27/DSqUdWJ7IeTgfc5mima4fLG6bDTrv6VzlmI27G/OGJsWrs/Sr+44
LqAir9WGjJx8zfD2M1oVrnZQGKdAIBLCGNqhhBIEG95YpLba3RtpJc088SOxVX0q8af7SzkNkd8n
u5B7Yb4VyZVmRARFEffZfnZRwki+MegKETXh33qkFPH0D9TCRxq7660uTffhbA6JjhlcIBlKZWFp
iNEh/6Y02hhi6BJ+LqvWOaDQcD8DzfZRlGnX36DbJbIgX74MKf7perJpWcqHXbv5M/M62zw1QDM7
j+u+y9AozcVRjW26yO1F8lH5lEzshCnxx9EQ/pUMszXRS5pF3NlTbwOGNnrgMNsLZbdL8SL0zTTm
FTGwuAiN1UYFDiUFKjHj72VI9kUR5V+8TAgZIbAtGFph80+0iMBwpEf39rO1lsDl5DuNYDXHsWyY
N0cDCNBLHHyMivOwVV1lByt/9J97o3D6zgPsh22ojQhp4fzSFRx0LA1uvjzVhP+YCTy/TP3QTIha
/BT/uxB2jarrA8cGgfqtG0doxP1ILpHwkh3Sm+Z9pQ+2+Fk5vKoTTpHMZwlqB3b/4ZkAgwbE+7bh
P9JnR/xXbBRybyGjgTgKZ2HgVMPgSa+WcD3S6aYxY/BuHauUR/vhT1V/0YDOr0kM/dgzmO61PX84
3me4yAfzRjRGm6MMTl7C9T0Vg4mW7YTSGsHc6u/cM6Bare4ISG8Ue//GHNT7hvc2APCg6PDoNa6g
xORsTcEeJjhyydsJYHCPKF7JCgTSPvVSbO7bYLe/Z2G+PslVp8Tyyqv0Y6bOcq7HJoq4o9lbQrxH
31/Gu0nWaME9fzYbKVrt/J1FU5LcPedy/BcSvKw3eIi0JD4YqITEd1hX2PgAe7t666I8kHgx6l9Q
B3W4mVEZ+y/p0UYjz0S72pZzRwoSgi6jB+2tMY1wwilzEoI6KWkqDCHfTroSlEm5QIRy+WfjkcQK
hHLyIqhhowprh35e+FGStozQp4fp45AFejG4vgHgFBNwGgWFdH56ZboS/tPYh4+D3FSRRFydOoHr
EBb6RFO25i4CJo9Er1PH0I1VwXMQn4FuiF08lpHIo0xFW21tk5Fj2OF853LmDDMNbnkBE3gmbbl8
sdcOZnxAumnl1pAgg3QvS+y49g7ZxRiCSa4Rhn+dJ64z/i4iTpzIqLZAVa3EQopv6GPkyNOmtiKt
HBaa6lGldY0SEWDBwdWg5LYkqGscEnJf+7dU9XeGHaGSwIW8O0o/ORFa2iwy24mRLLDU7aA4R3AK
eYpGOwq9h/og8Bh8QukpOe8a8SGF9oksUEuPyoqo+7XIFYbb9vwubLmvVYZeZFfE3iDvZl3REObf
GUF3Kl8rVlUARwiXBJizuTTCXumROG3VBLGzPO64kS8yDEbOz2zQ4Wo0eClEolQ1N9nHEF4KJiNc
Elpt2MTPhEbcxyFV/PD7OwA22eTDpVACPVIWkzhjgTYj4iXNO5dyJ338WDEJ8GrAfkc346QSfTeI
dp5HpHDhXi9uM6TPIIVNZS8rNvr2Bfcy3tB9iLAscIYrXPhDkbmSMoPDXB/UZYLzKh35e+4nX+Kh
JfRJ4rTOsF5hq6PNRPKeA/1WYm/JtQ3sJM5AOcuhRnAbdLqtSrIcCIaxgx7y2n5t23JrTy6h45jI
So/nesccMfdw594a6saMnxTNJbVTahzaclJ702DfO3RsdgrmqKLzSwFnHlrsxKoo7+Ztt3iDjLBO
TjjphBQacLcdBzgU5reZvgNg1ACdZM1b1fPgFaJbQcTCCCZBG/oDvchxfFDLbsiQuvOR7H2C/DpS
iJAXiUSdPiHnwqfW32hin0JBXuDNachN40ZpuCHFcgbCGapoEzKvU/w0L092fBMHNI8Jb3Uqh/ZV
XVzu+m+HWaW/QNoJWIzdrO3iyZ4W9c4uL8qknmCmQUSi4iDEJ0aqlys24tfVmvG0Tn9UIqgKkC3h
z5I/ahnRSLyf7wNqBcK65xUf188AHzlpztnYL8AbNbP0DPc7oYd87F50Jem/mUiIeLM93AV4lRJb
gKp3sFbvyEvWPDucwykLgPVqMoIGVgz1WJNJldlLI9DmEnOWfUNgSoupYDxWLFmg8JqTR1JJOKMR
Jrk4ILBg5IPOZAuLSV8iVJLEigdbkXa7UQLz64RsjML6mdC/GW08EC65YGxuiONSE+RQ68Ci372F
R/mwjV8rCGd+vidokJ6Kh0LxpNDAjnUjBBJY9d4IX8e13jQbLn4hmq+8d6bkXta0LR9kTV5sLLBV
xC+v6Jbq563ixAUGJCXpWFAiZkd6o//9zPJxhdCu/o86gdmF7Iuba6R3AKRHnhfslXXMlGg6EACQ
WC4VxUIHixOVp1wYJTO5+Ky9Xsb6woBZIjkKpzTO9YVa+PF+Df4jBitLgQ7MumqVtzkyVf0pRdFh
5iiYH4Q87ZC/7xwU/EC+Q0zBR5c7cQEQlzfpB+lIh30Jn2vBXpxKNyEuzsCluW8vIVVEfdG65OjG
nXb33AnpfnDypkrf4lKE3cTLgNc473Wb2pRsGDW6CVu+n7zajBUALZ7SL5A095L6CwLrWhXDZrXL
8+OzAmNLmyeJAScD84GYe7NNnqVJz6FmyVVYURHPDgP/WWEhaEsWhG8ICVHrCJs4X4iogsOlc5FS
kfKeHZcq03PCEimjkEiivFH2FnnM9FUjP2FpjuoPQC2LGLQbYPLNDS+yrR9kWgf5P7vIlVU/HbY3
uhB9g4CZhjiCh3VTRLV6Cw8/PgZj5NjE1DxW9fjEXdQHj98idTJMklmCTMPuCScXjTkLlkZb6FxJ
lHOVWLqSJFjMn2YIITpPPqJU1r1dO1//+d2+Co/aJLHBzE9A+QuZW0HP1vxS7NpkzwlU9+rW4RZD
2owSbfEngwhL2JOcrzN9HFTLlsk811e3rQuP4Wk/TS2RkQXRJ7buCXBXkQOGZIhJ91CyIVKPLT/D
okrfHV9WGqw/ehZWajnECgTgeYogQw4B+0FAgEiL/iZNq6XHbjdo91Nt/8ujgsApnz+XdODmNxsL
lGi5uT49DFeMf/9haNwohiUPHv8YHH8zr5UO8r/VGh996tTaR51bULczgB/s1LKd/dqCefrNptG6
6LA/Ea6Ox2OAMB5kc5mAEtN//0eyDmJVuJqjyj9cE2ue6jLiz2SVs8kANIzDOPXFwxTE4TZPOfh9
eClutdR0C3pTQFwRZJbXpjHxOP4nAA3kkPp1LRsUgAv0bx41hvxNjwHA1muc2Idf4Nh03Yi6wdOL
QvBxUDyGu7WahFhlqqrYfwh5A6WG+6Cb13xuF98O8qpPrEEYmKcHwukaCXmxLQNZbyofLvb/GjPk
W/kGak+HBhgE5O6T2qAtZJxySp6ranuVV0OrqfxbL1kWwo9hQBT3pWe3pf0HDdlBiw/FDk1RgbZw
0mDLkON0bIXrJMlgwTEQodYb9ivjALRt5wAKhIaMR6k7ZxQUCBSNQMMrUtSKKgiW5z2A8m1jTuhJ
JkNU8TWf/TtDYGN3x40kxG8fqzTWjEdaC311X2hBghy7Ra9se2BEETqalpd1kwmdRUbMymivW5qA
4TUewZfjkciZiszhm5OKKhF8IsIOBC8fNv9z3CSEG0wLC2JgdzOLtO4H3gR4mXgLAWD2Wsyca3CP
59dbJ49kCsXM048+sIJSTqAL6LlZNUIA4jEIjhfNy4KFL8OKhaaFXsiboVBRLqCcB7bbqZ1ihq2i
H/2a/bTebJekFPrEqWDcS7ct4gkJiParIwWIIb10W3yGqGClB/1eUe314JdWVoazW6+NtKFAXS9K
SCb5tSH5SpKNyUALeNlXVGQKgwVrFWCd+r4oUeqefwTFsway1QzxrWtqWpAJplLunwE+5t6eKLV6
mqe/TkUNEYOP24KTKJkVE0m4lOp8Hoa+7btZ1szLoeYvhgD4kzGwJv2JRnBBLVquHlqZ5si2ae5Y
ZOWpyKPDs3r35k1tLUsHFznG+oN4UsKEnZ5Vl4lh08D554GsEpg1/UTnO4XQVKSI9c8Mhn770fzb
4eby+ROTBkQ9aedONMiuberSVmo1azkuaYP0MsljDKhyL/+IFJF3sQxwod9owhIh11Ib1jmpqA4h
Ze9PpWWooyHR22p8P+kJtLd1BfOX88Wo328944yu1eJTpXA/FvBXobfngCwT+kPVRNfCHVhxpkG4
G2FWUMn746iFAgV/44Mm3trGldi+rs9NBJdWDWsWIx2+2JNlY0akgP9asnDPLSykLmjElGXofhte
ZTzLhWi2pMx9o0ajk679Ia8+1MjBqhcFYbd/9gwzhz6X8bTDsu6uQycdRCix5WoS5mabTo1uJtKv
cl/lq1zxO90QPNFurK7EtjynKcMqX/6/fXUcO3xhoKmpaWnGageImfWGWmTXsnJyn4QtioiDxltT
pXatRvP25c9Q+HprzaG5Xb70hc3jHIxiJP26h+8NPMpEPFB30OTo9UIGuwIW5nwEkI5wFvCw5cON
QHtXzXa4KhH9I6OTkwZX7KdCcZjC+nnrBNhFwpCGzrQKHTgRuZZDRzNRr3T2fIa2twIx2be5NZ6x
0mkO/4WaERDDBAgavT2rQ6fW+9+wI5FUkuYTjLxvn4ld/OXR5ObGD5qBVDXMYX/TG+9jR4HWHP3I
sbYEPvAfuI/+MhLyLFXgbTGV8kilffgIDsff92b6pBLlu1anUnAV54i1wPA1WlvVD2DmkaBOLQkh
IutqTgkr8+mbTmkQmTlwdTwoI8qGJnpcX9KfuI+CeHCT+syKoobZ7/MGCwddJ7gvAXE8iPg2cRC2
YzNTsUHAfgE+w9b1V5GNb1voehemjuMQAQkvXmGkCIsn81lW/nfVJPCj/h/iemUr7Ld6HhvaOqVm
9QJIQnHZQgS4qjAuEKN7TcK07EB8/QFrRbozMmS/e7yd/X65GphGsTLU8UzdLchMv3WAkGXEXmKo
weIEmvbcTMIeYtPLkpkGhJ8F5QLZAHRzzNjAAlHrvXjIDf6xXXNYIQYFWLxiSOx9SqmViJI2xiaz
/SkBOUiJMf1sgCc4ioEZXHXc2Rt80atml1pOaJrYITbEpM/MCBhlv+ENdIrFxu2FJY8JZjwZYWyu
CmWOz2lsVkkjn6wb3XDc+7pBSle6Pu0tOJ+f5IJwST9DS+lgIHlasmlZhmxYWGEOo9nU1qp4h7HC
TSMUFnmn2rLRAQOlJpSAIST0sesahqbECPtS9aDBfJ3Bq63Jd5eqKpwAkGZh9Sj90fvyoc+f7mfZ
P6/awCAHwVG9bjjRk3EDBkcvZwz1UOUk6NsaTbsul1Lu512d/vCBW8kHCAz32dMgKcfGliXgylkD
1a9+Uj3Esbk47OrWypMbD3ZRtKEbIPqrhLfpTV4waznS5qFRxlmrjbY9NdhVQr9GwuI+YNTepjoE
ROWZm8Hw8MnJ5TXG29xj0QVIgU872oA35AzN3NNi6Z5Hu8UIHl9sIx5AFC9PC/DK1GyTJ3W+IogH
lmRtoxzzxiGUI4RPwu/fmYR8LG1VpGK6pHKvJsS8nHdN7I1kO0yBzE6fl8miHAEBN5b7NlAw+P0Z
f4Omlro6vipfvrN9qONGMNonrkADrpyfexD4z07rHKnMENai0jM1yPYv/oVQUSACuQC3BYLz+aWr
COo0Zcz9buDtwddVU2nI1IDa0QHoN6kFYC+rgKXSp9wDLNrhE09n/XKzWupSztmegEzU/MLQ0Q+3
MSc+ugnOS8zPdu7zUChKMoW94e/oKQQpC1REFIdFBHtLBZV1N26qCgWrkieCtbQ7ANm8nb/BH4b1
FzgvmONd1nBPnDXaDMjTacS+eUHJskHF1gBaMfVckeQMSDkplNXxSyumo+JA17yBoEEuniJ0Kx9y
kxE7pTtpFw2YjEQzKDdqP4yvDtxApjoLR0PgSAvxZjI/FL++ijREZLp0sBMBvujAVCdG/8tmjru3
hXkbmZc4fieZ0VjDB5ccFvbp+doR4ZcUZhWFzbnjfxOi9RbNIXOxrdV1uQiHJ8S9dlc/D1FU79Ll
7XsL86QvqnploRUtEYetO9uyvVy9oujzpYkUpOuRz8QoLtAH0kCWaQERN28U0t5r0D1Vg47MM9M8
QSujAgQoTJST0H+Y9z1+ls4JQWy3Iw7fWC7Sfmdhv7WRxYQhZmz+qfotTuqRmyfutB0iTz9xNf7h
7h79UzZQnT8qgcqkjGIGuOFchTPaF2IN+LsryGoLnMGYyVHQUyFyNmnTpxKRCaedd4+q7K6UNy/B
IrDLf8jnHqYsx/gLS15EE91XbtkO3RwUcLSoZLxtHvPFwCjr12oV0x8LUj02ujrfq63Ro+1IdSbY
0FW1RRhMjeV/02ApKFcfkV8KmT+8+pcdgF0d9VlRUOQfRh955Rt50Js79jceQQH9g38+REcuPot3
6hAxdJ11NMo+OSuX4IKbL6bIYvNf1cNP2OhYGbc7OcWnn5X2pKMSAsvz1yzKJB6UqNlqaDS+6VCn
KQZ1BqJSUBbPJDxiALpCvkbv8lBLUjgov1US7z7M93tya5OKI9bq1ocn2EGkuiR4XvzT9V/p6Mbf
NCjQ6hx7H1QZFHistVmz99CEt32ZKHCbud22cqd6+v3C9nZLnFadm8+ZTqve0ZwX/NuDXaSiCPyP
am++1EaBX382YxXmCZyU0znAre9zkvhg16HAfPaF65gXjK4GCIdPqgZGnxV3jzb2FHX5o/61AvC4
q6qDZSzIIDGaNndczLF7hl45+4mN5Dhqf+QnSAYGzVhPg1IrjkKTIFZoBKa7urDa8Fv9qn3UOh09
YQRJrrFxKBpqgHKHSMmJTVoDxV5j5nMVqgLY05/KSQvq4xEW6X6ajiMvZB2L5d3o1Bcg6Tn5YHR4
t1q23rlWbpwhoroShwg9rjLd3scFRmJgSc704zQ9eiK9ujF0Ri/hQ6ADhH/l1cLvCV8+YNhYX+Jd
YPu4Vy8PrGAbLnCzWz3OAVjf0Gy98w7CRFUC5nr1Ojq4KpkDq1YUquCHbsQhg7e0bLyQ6j1R/IZt
q3o1ThLf6MCQFGxay5MBXxGIS2AMQuqwQsJnEsisPP0tu9h0+9gRQk+kg2z1jHbeCr6VlyZ35KC0
kgKMVceOOHcPIMQmWOBp+Itg7e2A6n0jFRm9QHaw1Vr1vxOQ2xolk7mjaHFsDLVF6w3e6Bul9fXa
mJYHshyFkQhnRk+PjubjdW07UqVOIOQLApU3cen3UyChblN8dQU5SvzkxeavJRw6/qbYJrUv04By
YNXfhCYXqUVqEcaNjz2RTmxYhsNJvXk1Bew/d/8UHEwbV/p7d+hC+RwwCiPkkxFrBixXrguntKWQ
li2QDjWYkPSq2xL78IW8Nfj/YkXniZBpgsqTTZu7nJifUtVrFG9+yzUzqDZOVfKiD5QXR2C0t1sm
5JPniUoHTlBOdVU43vvTt1vnG668udYt0LiqKUjiEjlnANtTaeElzjpivSxExzHpEG6hEcuRy6qU
8cqTCRKIAHuoTc+UB6T+N99q+KdCDlciTfSRd7nEeRb4h1oUS+JXEerf6eSMLd3qvGqjpHrCDhaM
+gZ/VEbslMrtVI6lj4JFLCS+PQl9z19aWwk9XsoBmieCnxyXtXzbxiwn+ibXM5q3h4oeQ8L4twde
357lJY61u9sEdVYOd0gAFEf5t4lXZ+9Og/F3CVJ/grVnCXxdMwH/BN7z45Oy8reDIrRchYRpKJJY
lb6WVcwKwdkrVM8VFyR0Pb2go7mkNwXqsfjflRQ+WyvlFlL1bg9Z9Ag4GqGE2BWLusKXcKn6aGo+
1NbKgbfR9hu/aAeH+5IwuBNmXVtLi2a+1gTtaMRYhlS8o5DgxNTFwafmqDXdWjcItTqzuzsM2qU6
aEqI4BYGQ3MLd8ZeCQ44P2YOPty9dM596L4JgYwWUTabnGlkNbgta8RtnX942X6g9ZsKc2er3pJn
VQu8IIRfjyTEKQ4nEsGfkrLsrUDdqNgrGtX4+6tm9cuhBePTxsd2kyw+9+qm7TKvwxCtPCJ1WjBA
Z8Vz9ItEhw9eUtUNY7IGLmuLj3GOjqmhNsQKifnFQ7sg3wzODh+rrtiHxqQM3FdG3fqqq64Sg+VQ
x36IlaxG+kqvFtb7YEu6NuMG/UyQjsEd7HyGeEzp7JEKjkzGRT0NjrlZva6WpOB1VXX+wh1YoFsX
V27y0GQCZ8GVYtRRANvO0wzS2WUe1CcnFkC+8ZvX0XIkyWY3nLTyeFia+54ifB/ANgx2hok+nKh5
WFSw+WQCnkX0nnrgWbSijmnHqB+i2UZ/yuCmT+TJzgYb5+zUWdaNbAk4Jsm5inaWj+WlU1zoorv4
02GzhwHGTPO2mqzJ+zsIAeLoEbYFPmSfsCHXsPnYfuWF8ShJJ86cp5FSrliRVZ/RjdICQ25NI5OY
yUMMKZGTN9gECFvWD7P5r8Jvq9Ni25YXlNZOYhGlnp/ZkmJ/27YGuj+YYJfj06IsMyy6+aVQRS3F
mRHePiwoFaALdCxFav+BPhT1WsipqfayHnHXaDyhGf01nL27R4hNv0cpxW36225oLsBgenUy8ebi
57Zx0STrLZBGjuy2fOlE6QPSBULQRduEKt0I/NX+ussi6lhvOb0vmZXXFDxthBDWO8ISIQPXno9B
fqFUwCpqT6bsy9ONsSFf6y2bE7TlbTNSWNZfYs+Nj4b3NxCnRXVM3It1bU9sjSo/+X2STle9B0z/
1AmbmqQ7aC0SzLcTZtmsslduX0gY86jxdH+GWzq0NSJL6aMxJNnEheq1EDPD8SNMTtKTEy0XDYHt
qx+dacO4jN5UZxqa2/xhHmnIr20W3s/hpjTX5EfESJda2DPSr5QALT3JOTpg3jgCpZqs1WoOc+Ua
U04xykmXhZucTqeK0lpZ5IKU4YOPauzy0inscEGxybg4cIJnFD8WXAHh0p0DMVj8g/Dvw7Uh1xRl
INxo6/DD1C3UoNuFHVSDx7ixVQKHGkWuGHD03tb1gBISB7zBH4BqoIJ9x4Q/qLOjxO9fuYBfjD7f
fzBSulIFaM6m93nL5MNVEAErqmJlmir/OSFsIQh4uiTDITR3Yq18y4q6X5IHIugxsHmZg7zXO/Hq
Pgu7TrwrIWmIOkvFPClDb27hMJSCOs4PN3joZh4m9wOfXLWir1Qan4OnW4zvb5BmHxOsXAPNgFiA
9Jad5JRZmTwkJ1ZHE6t4Ta5L6LhSbqhkxybiEaXtw1FBpzzfF5O4li2Rf3BTSBuIJT+xQH6dOob/
JD+MjAep9dGpZn9UVCwG0/eXtdbRPsXtyVvr/YMIs3+RcOJGpKJj3j3exE9x1LuNk+mV7upxZkho
bkUMsaCKtexugAEgKlqw97JBmz0MWarYYwRLyPROd8ZSwRrDAVVgawXHXufWazarDER8itql6MFO
5BkOekb/6ru6ordz7rOqTTDaS3yY7nyu1gYeJXqYNKNh11bBtEDFWhnUndWS9S+zrCcJb+lavNnR
hJphpTbKIqXJdsqpFG5DteVNS6R4N/0dqE9ho4UmlQhmGq0NkFE4W6Nh+AFBRNLhTt6evw1+YB13
L5WynohjOuDsDuo1VuIfkrMNhC0VCWYnu8rBlfpPupSH2ZV0JcKk9Y6Bdu+nBKcOktaqXNvOw5ro
9igpRcKcV2mEWgy2tMo+Z2sLB+Q8bJl2k1hgC9OhvnaIpOVT4n3dHxCVrUr7yLJ6EXyBmX6c9ld1
m/KCokIEOiKEUojqYPUVaMn9LFnJcZo1cyi1F0WjkcGfOzuPJAFG+mjtjWsMZoQLz/lVrELyaRa9
PaUq7ELclawjhqauyHw7k0euNvD8rjmj06mSu+qd/+U2OIda+VddGhyLWYOkidH9oIe0CWKe0pZW
LlhfV2Uuy0I/04Rans2wPeQcTlhXH5bXATilk5GqsL/GDWm1W8fahCjCycgUXbHao+0UPN4S0z3Z
n5yDVMwIgf0nOGbvKkPu6p6gzPYYqLFrb1JfES9M6OZWl++MrqmbLqCVvMS6AaYWCv+djIMT6d+k
t24Ff96R4Zg08Acjj82p7VBHDlhNPyEaztVij02uNwShkymsyCpXBJ4U0vYd2SZhkUvx0TYosa0U
B0yHvoD0qZvwM/8gJiI17qHQlw+xCxCU98oFYxgo0r8kAqtn8CS/lo2V8oUFAZqyJKXkG9Fbi1X3
xyDkuzW/ZwQHxj2B8HtB/k9cQ+rNpyuNWYGkf0ha9BQ7fS3zzpHax67ZqkowJ7q3XqA2J+pOe8Ts
RVPFVdLO6NSVW9pe9nxVtWTWdTWCDu+nMocwVYDkYM+eswYZByYqC/P84dCKzH4aF3PTM35VSBT0
r576BszFK0HD13+m70URhKkgG7rfQsIPt1OudhsTNMaoUYalYXjI+sgnYLAWJN99YkivzjEiR7Wi
l+YYpyVqjlBVDM9aQZSowBXJkbgLVsyIEF7WiEkXsTdd+JTF6phUnpr2Tqqusn5OGroPQC2f7XaJ
kHjpmOH+YzarEB6LmTzCe79o1i3vdTskENew22EfBans97mFQUZxqA48b6NyVIoBX7OeE7gGM15j
3pim3Cuy9eJSSnxdqFTOhUdLXXpRMYROSL3LCHlUvebqX1Kn45aLJFOu0Ze7d+4z6gXkyOLMh70s
eJUsWWg4G7i/8X3BKqqD0mRHc0NwLj9CqKynncK38QVSnEL8eOOWClgoCp43aclACL5jhKhu0XGT
vzhZ6HwP31Bvt3mOe748XaIDpzz0w64VdmoBkWsjLu8GsbMBM+HTVS7umRTgE8g8OnoteC51FsWT
Rh2OOGxab6G6lFnzDslDWrxVJoqV7aZMYdWTDGI/OlnPakOa2V98tUynszysw/9ZwDpDscr4B+6V
I592ixWuUj4pAYkf9RuqbS6x0+Wb6yTYPWzSJDPM1EuIWP+S6k5vrRbyRKNRKpN5y+DMqgKjAVe1
0QL/8xZdOmPFLYnE6mKNNpaKR38pq6RyHebF9yMaOc5JEFn1u/WA4Q17mP0nH1IQp8r/kZ72e83p
eAYG9kW/5QMeBszpxEsksq7tfM5d0PCaib9/G+vpbtAMQw2JWQ5woJ3Q4GBd2BX0FZMXjzE80lOq
m2S8UBFY7wYE7RqGFsqPjW3D7b/q3mlwR851BNWwEBUYid9bCFbaz11ZxR2MGkt+9a0g4sGiX6LE
FugUcMN7VNumYofT/Qqi1Y/yrTItFTgeoDl07xb6c/P5uRX8jMWBakZKfUf71OSPC2OhNNDIz0Y/
RdcCXYHMKpHJlwo2BDlHyQppugoO0uk2dSyjmnw3eRLb4OxFcThTyU2H7OnEgtJstAaRYBzIRgZV
w3p05pIdpfS6slfmFoonSkAOSTUwaNm2OGq+2WlHTX5Mi4KzGmeUqvUqjsY6q5kE1IPMU8v4oD1D
JA7PoPNXmdFq3QKlgMCstGKhPiOKZKzwfUPbBjQ6tKTs0BGnjzp7j1ZB4U1ZMZRoEdrxIJ9UqXJa
hljIGn3cyCtFrVQKfDUiXxSt5APXe3oO2nrwqfm6RKyell8mXpVwdxJzWA9CTvt/bZTwpykHpHLI
mI2uW4yMt7cR17cah5Zx8p610LDfMUvhGEBoqU5wUhfX1cyAyXCKfsm7jsbaR+alb1rT6X6dN5f3
/6hjCBB/v4PqZBKFPGkRhuWTcU2mxiCwI4QHANkEWxJUqkLFdt6D/Dm2GRUyKkYVatrKlUulZfV5
y/go9fhS5qbxvz2oG3OhGpwzS+emqY7NX1VqV7jU6BMcajxbxXtpQDYp7JAupvxu9W4r50DAxgK/
bAk7K4fJgQOoGJx/4DjcF0/2tGH2k5Nev2cciXlWYsqXUKRUiT9xtsUwWpL2dXwlPEZXCbby344A
6gW9u8T1oOpBVF7S4Ds2QMqY5s26NQEA5QCZDlv3QEQyfoDgV0y47gVl0KJi3uNDsn16A5sqFSLr
s7Kod6GFdNDWuLZ/bcorIeodFcB8ad4sd9WnRbGXsL1XrvWMSoUvSatgeB9JLhbY3QrU9MBlQqcA
Edmc/kJs5vlVz6b4Z5gnvGz3S15onuPgi3FpXC8APb1Lcq9qxNhumbVHhqm1xgleGJJJTXNBYCZy
p2r7d5K0JjMvex5Nk+j6w74YVbmWm4+CHJHHQ1c4y9trAV+ZpKJGWnFP7bZNpangF0bnw1BJwDvP
4dK4gpwKsVLcE+vffW857wONY0EEfOs7ZSX3IX6RVuX+z81H5EQMU83Ns6B6n37bzh7cOxd1U1Nw
yWeszk4AMrE3g3rjo12JKscVUMwsnvnbD97uVPXkVbU/ATmr7TxurpIPOCIsWyhwfX3qe4P9nJo3
T8goS9PXUDHXkDiCEk8wxBMcwo2f0j/QkE/bCH6tBmvc3iPIyA29g1bjupvAUKPqUF/s5/XIn34S
3KM0TDwEWuMj7DyfXFJSnwz/cn2dI4hqjXtdDR8r8B/07SiehOsFwQPZ0ILv5L4uvrBX3WuYkQif
yvChX491HhJRkdggDqD8gGoq+FHYokWX0irpi/xgYN/R9Eb9bL7er/UXPZnqqdTkhz14UCAPwC8l
FjmUBtJ7Q5RB10vZH6dcsBENn0fKgaDCDPwejlomeB0HkURhjFQGIGE2Yx95DnJ/eajeWD/3XpDK
jHvS+eTxIlXlg9yGyGmdqhyAdhtd/vpSPCo1KZIlzHw99tgXeyLBx9YxzGndL5K3OqKiFsoiWylp
tCq1EEtvB7KswFl6/7hI/Dm6yVb2jHUq8VAgracfE8SLqmNdb5BZCxdBNdrFqtTw3GGHBvMXN36j
uoX3ztrnPrYcGnbWt38uQ0rTBu7E6zRrhJLJrcj1eLs7/FVmtRNiYjI5NFlbKd4NSH1rW6O5k30v
KgWa9/v/C5ecGPACxgOyuV9RUN8FQAu7J5+QF+y3IP2FWjIlV6DYXRGkec9hmvF1ZjceulxqM089
eB5U9e6SRS5FtyCMXGlkaofGGxfNYtifXxgsgDSm226hXnAzFAtIoiPSPoL0mzTyOjw/9O0zjOph
2s+1r+ZLQ44U++HDhHgZ7p6ZQLtGRDxMYZddSoF5gUeYSi5JK0gyvZO5T5+3hjoEXfKxveFuc10P
FHqNnm4/bKwEcgrHNjPXstOOGgAMAhDSRLTJu+ldPPo9bWrWU2NHjrlVnxwFbu+Pdo9CBUPVQ9FM
vUTL/t2+RbA+ERLe1/WxKim3XcoO0LC2mYHipDG5epv65JKGhoqhcOnm9Unp96V0V96PxwRzj8+N
7ot+5oHcYdwJ5gifwhXYkX/bgam8kFK/fKyzXSKG9GfJbaaLwqXpu6bN/+69GoCVDAs0hAYDjL+S
XdV/kBJw0l0inSjoKQwFeCNVW4PsbCQIOjtbMD1CuQ4Gd9FyEFbGTBLY00VncOYqMYMFcKe9TNhy
P3a8+1wZhzEmlffiRKiOswxnp7EWounbH9hlRrACzzWo36bNJ/UAW6WkiniJ+qIA9EuX3WGzIcVE
2bAGKRwM6rW25+iaQBa0eHLvR06U9o2p3fF4/rEQVWwDmYVnFLFXbUxa82Av1MF8sFTMdKsDZhsH
2UasRGENb1R+7iNCwYKgl1eIWyunfe7g51KgJL3dR/v2ijBlk+LkG1FxtdjtC1HxQZs4sOOeWyxB
q1XvEnJ6pjBUzQ/Lflh2D+GzF9+FN7LJf9Y5pvo7Fj0WhRoWmVkw/rOH+SolX05zqNpmeuoWMSSB
8VqpcOV0FnQqswPhtjEBKIpNG+XQWAhGrcFdlYtgUXwNxFz6cw892spQqDIMUsEVdTUHdMxF9HZH
OibA2rF9LUxfVvSiDGlxKEE3omhGGmXKKyf910qEfacDBCCTGSeyC5yByKG7VMAub8jHJB6CtF6r
R2C2lu88AhPT+TBiCstQZu2EauQi5giCIDonuQXs2xbgwKZYjiSU06V9VSQMnuGgRBQG7D1Hc0pO
DKtvGiIw0Lb4EPNJGH7rer0Ba6eidc5Uj8XZhA8kBI0n+8E6JLvuvM92oIwdXRYF7CNWZx0vsvdb
PsLiu1sAIXDDIyR2fmnq1/l7F7T41wtcmSzOABPvOTUFMpu9opr3WYsTni+xOwiyRkt8MXD3ZS3w
bWnOTSOWI//1Y4iZFXcw0SzW6w8MciPiXjyIZdmHtRCVHMunWxA3IQxghjhaHtg2nz8zutVQj0K9
X7gnER/lE6QAsoRiEL5xEepXqZE3SAFbZNq7CIU9y4I9u+mGtVFDxwcRt1qa9iiSzoiVpb/qmxfz
aspDa+cKqjvFqRXiRD71yrI1j0vA4tOBIZc804RfGvjGYbTltWJm0+sBzp1lZu++Kbkr4K+F9GbQ
KJ+d6NcqAJ0jxh6+C2VocbxJZkA1KG8FdpIZzoXmJAXxK/2aW2Ng7TbOeUxmKv/fZ4aeZj24py8K
SIy+pPIQNPMPxlQcg5YkaXhGEGZEuO+g99N6TAq2utwPvH45oYlvQNH1G1vA2CJYIzSFPHcxfpXD
gCpBrZNnOYPQ00zZwYVGvzgtddubwvXneCcpuVnlMMDzpvMckSXIRoH4cVVeJzpvN9CJIJoQVjyE
k9wzYzCbzlPSEVlvFKUpzej/WsH9xcXX9gmISRIebNf39Wz9U/LNHHJs6ege6UdIXsNVbF07yFLm
Q7jnzhhple/ZV5+nn5lZEXKdYCOpvnm5ci3pChr97W7J1gh/wkrsd6+c+P5stsrmuWEKbrCrO0ku
ErRvmSxv3lASZ9RxmY3yOZyj9Ra36Imw7ZwPlccc4cz/FSLOphCxa3mNviMLn0W9Z6ap373yGHp+
CPtXvL4HmkfKqMqDjWPn7F/KJlyUUs4TIY5/99AjVElafVKs4ODicnBgvlaQgWK5E1E89D0qKqGH
HgID11XLtEufpvOmONKTOxsSdwLTs+b0R+lbuxVTO7lbxto8GA8Q84jPyLmk/TVOnvtxF24eaQ6H
0JUhwmS7FtzM5Be7+DTQmCJK7vFa0n+xMeewq6w/+EWTM5xQYbVNI1RZ/pqheiY3sSHuzWjoOGa7
wVT22DrdMh23G81DXzdh/S+MbNLiWPMe5tXn84FpfD3S73M+HXVvqp4+ND32MDKFxoz9KLKkmrSC
/Jkgw6uQhIiSXXpapRhM0hccRqFOHZ5vTSB2rjlEtFIV8FzT/kcIc5IaR3BuUBN6Ns4roDUycs21
I/o/++rCnhBEjrdfgJiEzF11fyBPhhYTnUcX+uuLqlL+JfQDKRwJxjfr6jqFD/2oNUwX3ZbKzs5V
Y2Vy+7nqviMS8MCkBTTzSZbKBndiArurEi2kPlTUHbfS3Ml5FfM39Xn5srwcB22fWN8A6lRbHbVZ
JZO0xXIPaOVvQjypLDWyaSvEfnHWFaxajYjRX9MvlTcrQd3IEGPx4tAgf92UMTB+rC4dtncrfss0
55ox9FbSPisd0t+tseFA8J6wd2xDuc7C6FrfMPYPQZyyweCFijiKc2+k8AB5Xh/b457UO9B0qjLi
SVv5Soz8W9GpzrWyyF7ZxUuFehTrvtf44kXlZXde+3BpGYO91272+0idUFnru0d8FZygOMeYDMYW
y5ca9Op/2xaOcsLz1QzG1PaQKNfvb4GHtmzK2XtdNbtKUx7bKy1JHGndeXsGFFi2tZQDKlrjQZlt
uwkjE+lJVUj+SyK8svEIOVgYV077RpIRJqNktG8f+TUv9nEQVr9OqDi92zd/lljz8CbjfEWJbx/t
hRzr35DOjCtJesg607K8aYzCWIcb3FiT67GqMmnyx+8GEgE1OVA+he/JST5LNZmE1wNEuKk6/eRl
XSX+XLn7Uxt6C5fxJyaGiFwALXL6vtCIPp9Kr2MSghjWI4yU6PCk/kK9/Tanbg5N+zZxIAEdX/Gk
xVVh8DLtBz7SZ0HBIJwHdBxfCaiR2pJVpaPrBV+VPQXB1FS8H7UAiIlQidGalqdeZRSeWub/p67B
vU2wlNciLFNzvtBzeQdnE2Hp2meRIgfNNv+JINSdi0c4E1AhiDQ/3Sas14Vzo3X/sYlcePWYLdqG
mXokyUcfwZDiX/rFw+CjxXSa4xYz75fVzyNObY3S91z+r2Wrjv/Aucbokz+KkeWiY6aVR/XlSo1Y
cm9dHxspgXiA+kWKk6gxWxOyZkgI+54FRB2fV8WE6Gk1ls6pEWajpamCzak7aS1ihJ6mfgYdwA3C
SHbtkaf693a92HVEpG0Wiyg6bc0D1H9rI7md1G4Z3X8AHd8KFqANoX8rsRNxCKCxmhoGeHwJaGvr
bnOA4Doe8Gxc4Vnm160cHC9aa600UjKf1QfDoqxineuabqehtgKpr8rknk9FAjuZvonV8Pf8GvC+
HlWhpUhWPd9Fc18G2duf3uSn2/yV7INCAqLB74liBrdAYkxAYd2UhWB6ePLfFeH0jINpef4BA2fB
9ki/UaE4XGLt0cO9i+dbfq1ajNNrbolDuCwUCTVszHyZC7Y03OkpqobL1LwqjagZbZ1SDm/Vh8fr
eJD9bMYxSXrbn9DeeAAVoOTwq19PoUK+ttNofx0iwr/2aQpcaAKEUQHfZHw8j2Ai1Mruy2NAPdb9
LYfRzaPSONWOnj3hn7k3amSebWFyRnSFuxbXEPoLNayZJ4yL9l/AYXhfc8uzHOs2yKy75eWkFU3j
SKr0qAQA+P60otp0JEY+rVyRKOdmzAEqkYmwrHsZ0UxZYikS0zW7eTe4oUv5YuO8pIC4C26T3hVR
JWq0iDbVcyXu3NN0elCuVFCrBKSmAcDHhkeIEItimgmF90iDh5mzLDj3NQqMltspObE/3qdYB+F6
LvJ3LPav8E7B4YyPxgVny0NVcHbcwSDMV2KNWQEpwT7Aueh7WirRC0HvUXPRcUwKeTpPIjv7iJWe
/HRg3e3VafBq4I90OdkoYPPtFmSYmdEDqIqsKplrtrxg2p5uSXu4X2OjJao/hkFkl8ylUuxmK+It
y/DxjPInb8+KSo0af3npN59BlnJDPHvvq/E2Hk8QbUN+/bzqVsRU80+sxYWFR2VD+Mzcz7pUVHF9
C9uoTV1ETrddjg0nBZNRb+6mbnVqDyHXLbhWo7jEwgf4nSAQ9GerPqoZoCCWDd7s5Y9jOainazTS
L6pi12qtf+WQeRBFUGjChi46CFsn2ocuYn8TUNc9PeqDPQoWm0ye9uLc43xVwMoJ9Isfj7/STP+q
nsrizcVGSYVlpuD9NgYIT5xZpenLi16XMYsJJ5w7NqU/ztzVFCWAsEw5CxdZUf5HopYk+C47V4rm
axTTv1WwiiNSTrefPfaK+Y2DhfJ6FnWQ+6vAF1RV7emKkKIl23C0NYOXDwFHcpLhg7tNNs6pTbtP
xcrS71qrV182RIAuH/svSxZoYBOpB0LPKNFpd43pm+rU4lUuHyvHbBOhCOf9t68Pbk5EgxBKi8yr
j2YHOyZTlbjIGTz4u6AnfZn20S/0WNXtfSyefTyUAcXVYSLR1xr0jd7dlEJfrVcxDbSH3N69WXVF
7OkNZwPUnX8hh73PB4GvsfE4VrUFvpLGZSo1M9uFnrI/2tmcwSfObQiJiblf+OvjITAuE5vnG7KK
5ezfs3jsYufCETpl5PuKunAzkPt086svZOcCRRQsndhA/V+9xyynDC7Uni5An/3eeVaPtEdpS29j
JRce4/Kds2uXj4/tmbbMUuZZHg+kRy6NhPFyFLWmGS8uhNvGmT63m3wHBMaaj7fXWXpqqh0YvXwp
vKuzJtIuzhXDokRKxbrdzatpTpZEzpvF5lOLrR4CZ8Dlj2cfb2PM0CbvPM+Dz3NTCMdFta3GrLuo
Vwt9A3uHwsCLC5ie2Pukyd18kUp+1YmzIxC8mMMheBmqS2sWxmxnL9GoLPIK8nxn3f6fZaG5zdeh
0PuUC35oHhqkhhwyX585m6ImumNmnjbBQbY5WE3BOKzjX5AC88/wpt4QPuYmz5MFdKHVLQPpkqvD
dVkiMGFejjooAGUox0rSc7GhA7bQVhPOihThyZom+KAnGZlsY/TQDpEAM92blJ+99FamBlhbgnpc
IgjnwFKuKKYD8guBsY60V4Xf8MkUhBZKmGUfEVvCKwhUea42xu0SM4WnAns6J+GcB2bYqlEHTnpd
eDPz5mxymgqXmlhRJyBq9qf2gBYM2FM9IPyrsaXuZS1W/K47hUmlnLBPKBh3V2WMDvT8GTuFxjTt
9sHOaYt9Tuym03Mgs8yOOjmRBJuF2ahm7oZH8r/TmEU1pNCoC6QQUD45h4hPh7PRor4R0rJ/G68R
v5H11rGI7W6g8At5poSrUa4za79KYWAohtpGVwwP6CXxRSpdlIpvK2OtjhlR3es34veI/T6FO9qY
aS5KjCW4JZ93LS3lAmTJgRtDCq8tk22WUM5aBrnATIkRSmEkNQAxDLBIKqb5xHXy8Kmhxvf66Uld
ioYIlEvR3rSIf0aEkTIqZRx4QNTRVS/oD567PquNPDW1OTyBheyQzOm1T8YjHwBvj2/4Cicvt1wI
mY4rkWsROzeJ7s9hymCn5qn/k9fGJeR01cyoirZxr4ktXHU7JJp3deHSZ/3TDDq74rXEaIJ4lk1y
s3ZbI71QvY0jMaZ1X1I6L5b/bbiHzMPv0dEjxyikVncS6m7fb/OD0Y/YWRMwUm50CVCnv2PybR0E
bMyWynSzCe9bs8fT9d48YLaLTM7AIv1XcNQ4SXxKmFAljNqdfNoMPLin3sitHA84GJKFaHcyPfHQ
eDVxIKN93zZhwtt3hMdC2YJbomTkQZPfD1+dMt5r1HkqYWT4+hFr0ErMMISbp6BKQ9Ws1CZL0K/I
Vjj6dtsfRwZ2JgXYKxL4JpSvxt3F/7gHuqxMupx5vB3U7DLj8DpcR/1to4FAf0Adzu00pYeCwivX
K8ycAY7R5lDUBk4oMad0aWLBiGsFCXl09zmLWs4RQHdRLOJzhCtKUlSo7upZ3ydCmqkPfDbPF90n
CYFsRYy+Yd4BXZv4/y9pUgZAyIzh48Rq/SNltsVEQHmZzJKgYImXqXPjfkQixT9w3UaZfhay/vzA
sHMAZ7vXBYfwVOPoIWy8CK07hNvek6346Kc0lJ7JZAkRsQUgRIip6GI5HomejzTLGlcO7AJhaAu1
0nY1F2wXOpU3aLOjD3XXHYccvJkhFZlfW+gPfjZyEJsz8K+G6/qlJCPf7sQB8PwUdhj9nolmpO/v
oTUFO8bcxR+6RqBJVySZSHlHnagcYV4c2LeUZHo+eRiPIT83OS7bLzLq5qr6ImvhtEWLWxPLL4X6
b0aaVZEUBel2cE6R+wrGZ8brzHzBPKGQvoDlS1zyNIGFLeygrvUr9yj/U6osUTwxLuxW37Q7cOgS
SRuvCMr5/Rk5O4uqlSg9lAj3WAB4QFyzvTe2k1CMz9kV+0RDiaipNMtUHJBz2zUiqgZCOINbLsqy
EGofghHiSJBTkRaOeTcJWLNeItD1W1H5EwbXpVDWVqi7II620xZ/7bg3BcpkRvrnNf0YZfHRFyYU
zdSLdsZkAVsv8HwhB9mZu3y1t+YMZXSS7sXqUGdi9f4TpWaY+DJnkxDu6tXUjnl7mOPk13jRuNyL
1rs/dIknmppPD3sroIRLF98eesPuprBjQEKari+br6shzarO0XLaWSEXcq9v8A+WPmYLLhMT5s2m
MERWxaLokjEyNWH0WwwOsyw3Zj/gFsv0KbpLJLhzQQ/s4t8AucENCuQmSyJJQJNNmo9hg7cnUe1G
Lo16TuJmcrLzP1f9h/W41eWyRYRl32Zs6rEDqtg+9I5gwuJtbaw3gAvsn7qdVC7kaz6QYEQhw3Cp
utCLv1A8TxO/N0fpQOFS8uqtZagDDyzk96X3FpIB/vo42Jv1eLZso2qOTRgbpNc97h869T1jF3Xf
fU8Bb5jilGcqIFQlQIN8L6B4AwKaeRw7EvnHr1U7T649IZrPxcXH5nJ2qo6AXThSg2EjxkXJt3+f
tegsr8ssVqYleDym/xZiqdwDR1Fz92FlDJDq8V4ysGmoBZ+/1/nI6XgsLZiQylrELLu2VWJuRtWm
DTgGhvZRJOT3Ni4hzr4hTn7UwZSwS71GG06Wcdz/tU6sRSeg8rBWEwltYEXW5pV2eYPVfv4VzlsG
yBwGdm6xJ21s5WMK4cnqmi6KJjNQl8WjyGr42b85Z3YzJnJOHI8REFNruYufSybhoWtaHoJDQ8lg
tRvWOl+jzoJSLGKpJvwyayxy+cOBswRU4cl41KdVWTLRUMEGz8dULdMWUNaMjufr2CNQnjYLsiNe
IIyndHiTuWoUBSnehbmCepEc2gKa9Q+t3mU4Mw0yL4lWJhioL+KhfREwYpGOMq6RUEMdcBFldGor
IiDJppFlJNVKq4GicTTiyOtwhwzXOtlv3G9S/XISaEYwajVhDbFtEstEQv+VL5uHczuiAkG+QR9J
POEgECQ4SuK1d3yo4NDijN5rrQ1PBnpbmkcdJgGI7Os6nK16yAWBzsUBBkR3nRBr8TiTS2I1aRaD
ozJwN3NNx5aig4pP7lf6INBY+cNeByV22o3D8qgGawKG7lsjMhtoup2quoQt2fDJ3ModAk2Ngg4f
m0LodPhYhjfcVgPN+4HJNQFyHlYOE2DB9w8D9dwzvOroUZrg3TJOiI7nECbuQS28DFV4nWt40MZi
VfYpZlhSE95o2ZAP6ud+hGVqj5UKpTFReJv503hLUNq7QaLP1tGHuRn9oDhiH6SGU6iZj9FNHKXE
R8R/GPpkIBO2xF5GX3iiA9lK/HD5B8lie1OSVm5EVEK41ffhNWMX0igWF1aSxrLyrFhZoFEKuYw3
a+Jxe302eGCtfYMSDSzGjYAzZX7GXpCu3RrB9nJVfkpjBNCK8/ftbV4AWiREpnxtYKdswFyy31eQ
5YM34KND66OhhIXlIZAIIMjv3b4+572/OlzYKHlwMbbhXiK6Telfr+sw/1hBm/rx2Mcr+e/KjqH+
1MAd0yRMV7iipk2iicUVE0Ez9WBzLEdFHnGD7EqGze+dAIx8MW29R5DGiJMQlCt4rY2xhATa/Tqo
pcDMHurTU4VAeonj8KR2olXES5i4OMiiSKQWNcin1srqRVs2aOkGOgs4S1fgt4OTrX8Obel2Ff7a
wVuqHpIZ9FoATcRf9eM/gmdZzqdXDBYRvNOI89sTP5pn5wXbC1Edz5fccmu3B4d8NHfYFrwZHrvH
LLGc1rfmpeukJhzyZY/sXvoANUJ/t4MKvK1W0v4Yg7wpAOpZMfX6iKkgUBUfdqeWUtfU0dUvml9n
4yBj+URc/4iHGUGgQEkguq2dxZR+LvP9EoHdBxaTS/C1BJ6KTE/7o66c8yG5/h4=
`protect end_protected
